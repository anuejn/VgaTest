library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity picture is
	port (
		vState : in std_logic_vector(15 downto 0);
		hState : in std_logic_vector(15 downto 0);
		r : out std_logic;
		g : out std_logic;
		b : out std_logic
	);
end entity picture;

architecture first of picture is
	
begin
	r <= '1' when vState < 100 else '0';
	g <= '1' when hState > 300 else '0';
	b <= '1' when vState * vState < 300*400 else '0';
	
end architecture first;

architecture me of picture is
	signal rgb : std_logic_vector(2 downto 0);
	
begin
	r <= rgb(0);
	g <= rgb(1);
	b <= rgb(2);
	
	rgb <= (others => '1') when ((vState = 0) and (hState = 589)) or
								((vState = 0) and (hState = 590)) or
								((vState = 0) and (hState = 591)) or
								((vState = 0) and (hState = 592)) or
								((vState = 0) and (hState = 593)) or
								((vState = 0) and (hState = 594)) or
								((vState = 0) and (hState = 595)) or
								((vState = 0) and (hState = 596)) or
								((vState = 0) and (hState = 597)) or
								((vState = 0) and (hState = 598)) or
								((vState = 1) and (hState = 590)) or
								((vState = 1) and (hState = 591)) or
								((vState = 1) and (hState = 592)) or
								((vState = 1) and (hState = 593)) or
								((vState = 1) and (hState = 594)) or
								((vState = 1) and (hState = 595)) or
								((vState = 1) and (hState = 596)) or
								((vState = 1) and (hState = 597)) or
								((vState = 1) and (hState = 598)) or
								((vState = 1) and (hState = 599)) or
								((vState = 2) and (hState = 591)) or
								((vState = 2) and (hState = 592)) or
								((vState = 2) and (hState = 593)) or
								((vState = 2) and (hState = 597)) or
								((vState = 2) and (hState = 598)) or
								((vState = 2) and (hState = 599)) or
								((vState = 3) and (hState = 593)) or
								((vState = 3) and (hState = 594)) or
								((vState = 3) and (hState = 595)) or
								((vState = 3) and (hState = 596)) or
								((vState = 3) and (hState = 597)) or
								((vState = 3) and (hState = 598)) or
								((vState = 3) and (hState = 599)) or
								((vState = 4) and (hState = 594)) or
								((vState = 4) and (hState = 595)) or
								((vState = 4) and (hState = 596)) or
								((vState = 4) and (hState = 597)) or
								((vState = 5) and (hState = 593)) or
								((vState = 5) and (hState = 594)) or
								((vState = 5) and (hState = 595)) or
								((vState = 5) and (hState = 596)) or
								((vState = 5) and (hState = 597)) or
								((vState = 6) and (hState = 591)) or
								((vState = 6) and (hState = 592)) or
								((vState = 6) and (hState = 593)) or
								((vState = 6) and (hState = 596)) or
								((vState = 6) and (hState = 597)) or
								((vState = 6) and (hState = 598)) or
								((vState = 7) and (hState = 590)) or
								((vState = 7) and (hState = 591)) or
								((vState = 7) and (hState = 592)) or
								((vState = 7) and (hState = 596)) or
								((vState = 7) and (hState = 597)) or
								((vState = 8) and (hState = 588)) or
								((vState = 8) and (hState = 589)) or
								((vState = 8) and (hState = 590)) or
								((vState = 8) and (hState = 591)) or
								((vState = 8) and (hState = 595)) or
								((vState = 8) and (hState = 596)) or
								((vState = 9) and (hState = 587)) or
								((vState = 9) and (hState = 588)) or
								((vState = 9) and (hState = 589)) or
								((vState = 9) and (hState = 590)) or
								((vState = 9) and (hState = 594)) or
								((vState = 9) and (hState = 595)) or
								((vState = 10) and (hState = 587)) or
								((vState = 10) and (hState = 588)) or
								((vState = 10) and (hState = 589)) or
								((vState = 10) and (hState = 590)) or
								((vState = 10) and (hState = 593)) or
								((vState = 10) and (hState = 594)) or
								((vState = 10) and (hState = 595)) or
								((vState = 11) and (hState = 578)) or
								((vState = 11) and (hState = 579)) or
								((vState = 11) and (hState = 582)) or
								((vState = 11) and (hState = 583)) or
								((vState = 11) and (hState = 587)) or
								((vState = 11) and (hState = 588)) or
								((vState = 11) and (hState = 593)) or
								((vState = 11) and (hState = 594)) or
								((vState = 12) and (hState = 579)) or
								((vState = 12) and (hState = 580)) or
								((vState = 12) and (hState = 581)) or
								((vState = 12) and (hState = 582)) or
								((vState = 12) and (hState = 583)) or
								((vState = 12) and (hState = 584)) or
								((vState = 12) and (hState = 585)) or
								((vState = 12) and (hState = 586)) or
								((vState = 12) and (hState = 587)) or
								((vState = 12) and (hState = 592)) or
								((vState = 12) and (hState = 593)) or
								((vState = 13) and (hState = 579)) or
								((vState = 13) and (hState = 580)) or
								((vState = 13) and (hState = 581)) or
								((vState = 13) and (hState = 582)) or
								((vState = 13) and (hState = 584)) or
								((vState = 13) and (hState = 585)) or
								((vState = 13) and (hState = 586)) or
								((vState = 13) and (hState = 591)) or
								((vState = 13) and (hState = 592)) or
								((vState = 14) and (hState = 577)) or
								((vState = 14) and (hState = 578)) or
								((vState = 14) and (hState = 579)) or
								((vState = 14) and (hState = 580)) or
								((vState = 14) and (hState = 581)) or
								((vState = 14) and (hState = 582)) or
								((vState = 14) and (hState = 583)) or
								((vState = 14) and (hState = 584)) or
								((vState = 14) and (hState = 585)) or
								((vState = 14) and (hState = 586)) or
								((vState = 14) and (hState = 590)) or
								((vState = 14) and (hState = 591)) or
								((vState = 14) and (hState = 592)) or
								((vState = 14) and (hState = 594)) or
								((vState = 14) and (hState = 595)) or
								((vState = 14) and (hState = 596)) or
								((vState = 14) and (hState = 597)) or
								((vState = 15) and (hState = 576)) or
								((vState = 15) and (hState = 577)) or
								((vState = 15) and (hState = 578)) or
								((vState = 15) and (hState = 579)) or
								((vState = 15) and (hState = 580)) or
								((vState = 15) and (hState = 581)) or
								((vState = 15) and (hState = 582)) or
								((vState = 15) and (hState = 583)) or
								((vState = 15) and (hState = 584)) or
								((vState = 15) and (hState = 585)) or
								((vState = 15) and (hState = 586)) or
								((vState = 15) and (hState = 587)) or
								((vState = 15) and (hState = 589)) or
								((vState = 15) and (hState = 590)) or
								((vState = 15) and (hState = 591)) or
								((vState = 15) and (hState = 592)) or
								((vState = 15) and (hState = 593)) or
								((vState = 15) and (hState = 594)) or
								((vState = 15) and (hState = 595)) or
								((vState = 15) and (hState = 596)) or
								((vState = 15) and (hState = 597)) or
								((vState = 16) and (hState = 574)) or
								((vState = 16) and (hState = 575)) or
								((vState = 16) and (hState = 576)) or
								((vState = 16) and (hState = 577)) or
								((vState = 16) and (hState = 579)) or
								((vState = 16) and (hState = 580)) or
								((vState = 16) and (hState = 581)) or
								((vState = 16) and (hState = 582)) or
								((vState = 16) and (hState = 583)) or
								((vState = 16) and (hState = 584)) or
								((vState = 16) and (hState = 585)) or
								((vState = 16) and (hState = 586)) or
								((vState = 16) and (hState = 587)) or
								((vState = 16) and (hState = 588)) or
								((vState = 16) and (hState = 589)) or
								((vState = 16) and (hState = 590)) or
								((vState = 16) and (hState = 591)) or
								((vState = 16) and (hState = 592)) or
								((vState = 16) and (hState = 593)) or
								((vState = 16) and (hState = 594)) or
								((vState = 16) and (hState = 595)) or
								((vState = 17) and (hState = 574)) or
								((vState = 17) and (hState = 575)) or
								((vState = 17) and (hState = 576)) or
								((vState = 17) and (hState = 580)) or
								((vState = 17) and (hState = 581)) or
								((vState = 17) and (hState = 582)) or
								((vState = 17) and (hState = 583)) or
								((vState = 17) and (hState = 584)) or
								((vState = 17) and (hState = 585)) or
								((vState = 17) and (hState = 586)) or
								((vState = 17) and (hState = 587)) or
								((vState = 17) and (hState = 588)) or
								((vState = 17) and (hState = 589)) or
								((vState = 17) and (hState = 590)) or
								((vState = 17) and (hState = 592)) or
								((vState = 17) and (hState = 593)) or
								((vState = 17) and (hState = 594)) or
								((vState = 18) and (hState = 572)) or
								((vState = 18) and (hState = 573)) or
								((vState = 18) and (hState = 574)) or
								((vState = 18) and (hState = 575)) or
								((vState = 18) and (hState = 583)) or
								((vState = 18) and (hState = 584)) or
								((vState = 18) and (hState = 585)) or
								((vState = 18) and (hState = 586)) or
								((vState = 18) and (hState = 587)) or
								((vState = 18) and (hState = 588)) or
								((vState = 18) and (hState = 589)) or
								((vState = 18) and (hState = 592)) or
								((vState = 18) and (hState = 593)) or
								((vState = 18) and (hState = 594)) or
								((vState = 19) and (hState = 571)) or
								((vState = 19) and (hState = 572)) or
								((vState = 19) and (hState = 573)) or
								((vState = 19) and (hState = 584)) or
								((vState = 19) and (hState = 585)) or
								((vState = 19) and (hState = 586)) or
								((vState = 19) and (hState = 587)) or
								((vState = 19) and (hState = 588)) or
								((vState = 19) and (hState = 589)) or
								((vState = 19) and (hState = 593)) or
								((vState = 19) and (hState = 594)) or
								((vState = 20) and (hState = 571)) or
								((vState = 20) and (hState = 572)) or
								((vState = 20) and (hState = 585)) or
								((vState = 20) and (hState = 586)) or
								((vState = 20) and (hState = 587)) or
								((vState = 20) and (hState = 588)) or
								((vState = 20) and (hState = 589)) or
								((vState = 20) and (hState = 590)) or
								((vState = 20) and (hState = 593)) or
								((vState = 20) and (hState = 594)) or
								((vState = 21) and (hState = 585)) or
								((vState = 21) and (hState = 586)) or
								((vState = 21) and (hState = 587)) or
								((vState = 21) and (hState = 588)) or
								((vState = 21) and (hState = 589)) or
								((vState = 21) and (hState = 590)) or
								((vState = 21) and (hState = 591)) or
								((vState = 21) and (hState = 593)) or
								((vState = 21) and (hState = 594)) or
								((vState = 21) and (hState = 595)) or
								((vState = 21) and (hState = 596)) or
								((vState = 21) and (hState = 597)) or
								((vState = 21) and (hState = 598)) or
								((vState = 21) and (hState = 599)) or
								((vState = 22) and (hState = 584)) or
								((vState = 22) and (hState = 585)) or
								((vState = 22) and (hState = 586)) or
								((vState = 22) and (hState = 587)) or
								((vState = 22) and (hState = 588)) or
								((vState = 22) and (hState = 589)) or
								((vState = 22) and (hState = 590)) or
								((vState = 22) and (hState = 591)) or
								((vState = 22) and (hState = 592)) or
								((vState = 22) and (hState = 593)) or
								((vState = 22) and (hState = 594)) or
								((vState = 22) and (hState = 595)) or
								((vState = 22) and (hState = 596)) or
								((vState = 22) and (hState = 597)) or
								((vState = 22) and (hState = 598)) or
								((vState = 22) and (hState = 599)) or
								((vState = 23) and (hState = 578)) or
								((vState = 23) and (hState = 579)) or
								((vState = 23) and (hState = 580)) or
								((vState = 23) and (hState = 581)) or
								((vState = 23) and (hState = 582)) or
								((vState = 23) and (hState = 583)) or
								((vState = 23) and (hState = 584)) or
								((vState = 23) and (hState = 585)) or
								((vState = 23) and (hState = 586)) or
								((vState = 23) and (hState = 587)) or
								((vState = 23) and (hState = 588)) or
								((vState = 23) and (hState = 589)) or
								((vState = 23) and (hState = 590)) or
								((vState = 23) and (hState = 591)) or
								((vState = 23) and (hState = 592)) or
								((vState = 23) and (hState = 593)) or
								((vState = 23) and (hState = 594)) or
								((vState = 23) and (hState = 595)) or
								((vState = 24) and (hState = 572)) or
								((vState = 24) and (hState = 573)) or
								((vState = 24) and (hState = 574)) or
								((vState = 24) and (hState = 575)) or
								((vState = 24) and (hState = 576)) or
								((vState = 24) and (hState = 577)) or
								((vState = 24) and (hState = 578)) or
								((vState = 24) and (hState = 579)) or
								((vState = 24) and (hState = 580)) or
								((vState = 24) and (hState = 581)) or
								((vState = 24) and (hState = 582)) or
								((vState = 24) and (hState = 583)) or
								((vState = 24) and (hState = 584)) or
								((vState = 24) and (hState = 585)) or
								((vState = 24) and (hState = 586)) or
								((vState = 24) and (hState = 587)) or
								((vState = 24) and (hState = 588)) or
								((vState = 24) and (hState = 589)) or
								((vState = 24) and (hState = 590)) or
								((vState = 24) and (hState = 591)) or
								((vState = 24) and (hState = 592)) or
								((vState = 24) and (hState = 593)) or
								((vState = 24) and (hState = 594)) or
								((vState = 24) and (hState = 595)) or
								((vState = 24) and (hState = 596)) or
								((vState = 24) and (hState = 597)) or
								((vState = 25) and (hState = 572)) or
								((vState = 25) and (hState = 573)) or
								((vState = 25) and (hState = 574)) or
								((vState = 25) and (hState = 575)) or
								((vState = 25) and (hState = 576)) or
								((vState = 25) and (hState = 577)) or
								((vState = 25) and (hState = 578)) or
								((vState = 25) and (hState = 581)) or
								((vState = 25) and (hState = 582)) or
								((vState = 25) and (hState = 583)) or
								((vState = 25) and (hState = 585)) or
								((vState = 25) and (hState = 586)) or
								((vState = 25) and (hState = 588)) or
								((vState = 25) and (hState = 589)) or
								((vState = 25) and (hState = 592)) or
								((vState = 25) and (hState = 593)) or
								((vState = 25) and (hState = 594)) or
								((vState = 25) and (hState = 595)) or
								((vState = 25) and (hState = 596)) or
								((vState = 25) and (hState = 597)) or
								((vState = 25) and (hState = 598)) or
								((vState = 26) and (hState = 503)) or
								((vState = 26) and (hState = 504)) or
								((vState = 26) and (hState = 505)) or
								((vState = 26) and (hState = 571)) or
								((vState = 26) and (hState = 572)) or
								((vState = 26) and (hState = 573)) or
								((vState = 26) and (hState = 576)) or
								((vState = 26) and (hState = 577)) or
								((vState = 26) and (hState = 580)) or
								((vState = 26) and (hState = 581)) or
								((vState = 26) and (hState = 582)) or
								((vState = 26) and (hState = 585)) or
								((vState = 26) and (hState = 586)) or
								((vState = 26) and (hState = 587)) or
								((vState = 26) and (hState = 588)) or
								((vState = 26) and (hState = 593)) or
								((vState = 26) and (hState = 594)) or
								((vState = 26) and (hState = 595)) or
								((vState = 26) and (hState = 596)) or
								((vState = 26) and (hState = 598)) or
								((vState = 26) and (hState = 599)) or
								((vState = 27) and (hState = 495)) or
								((vState = 27) and (hState = 496)) or
								((vState = 27) and (hState = 497)) or
								((vState = 27) and (hState = 501)) or
								((vState = 27) and (hState = 502)) or
								((vState = 27) and (hState = 503)) or
								((vState = 27) and (hState = 504)) or
								((vState = 27) and (hState = 571)) or
								((vState = 27) and (hState = 572)) or
								((vState = 27) and (hState = 576)) or
								((vState = 27) and (hState = 577)) or
								((vState = 27) and (hState = 580)) or
								((vState = 27) and (hState = 581)) or
								((vState = 27) and (hState = 584)) or
								((vState = 27) and (hState = 585)) or
								((vState = 27) and (hState = 586)) or
								((vState = 27) and (hState = 587)) or
								((vState = 27) and (hState = 588)) or
								((vState = 27) and (hState = 594)) or
								((vState = 27) and (hState = 595)) or
								((vState = 27) and (hState = 596)) or
								((vState = 28) and (hState = 491)) or
								((vState = 28) and (hState = 492)) or
								((vState = 28) and (hState = 493)) or
								((vState = 28) and (hState = 494)) or
								((vState = 28) and (hState = 495)) or
								((vState = 28) and (hState = 496)) or
								((vState = 28) and (hState = 497)) or
								((vState = 28) and (hState = 498)) or
								((vState = 28) and (hState = 499)) or
								((vState = 28) and (hState = 500)) or
								((vState = 28) and (hState = 501)) or
								((vState = 28) and (hState = 502)) or
								((vState = 28) and (hState = 503)) or
								((vState = 28) and (hState = 572)) or
								((vState = 28) and (hState = 576)) or
								((vState = 28) and (hState = 577)) or
								((vState = 28) and (hState = 579)) or
								((vState = 28) and (hState = 580)) or
								((vState = 28) and (hState = 584)) or
								((vState = 28) and (hState = 585)) or
								((vState = 28) and (hState = 586)) or
								((vState = 28) and (hState = 587)) or
								((vState = 28) and (hState = 588)) or
								((vState = 28) and (hState = 595)) or
								((vState = 28) and (hState = 596)) or
								((vState = 29) and (hState = 486)) or
								((vState = 29) and (hState = 487)) or
								((vState = 29) and (hState = 488)) or
								((vState = 29) and (hState = 489)) or
								((vState = 29) and (hState = 490)) or
								((vState = 29) and (hState = 491)) or
								((vState = 29) and (hState = 492)) or
								((vState = 29) and (hState = 493)) or
								((vState = 29) and (hState = 494)) or
								((vState = 29) and (hState = 498)) or
								((vState = 29) and (hState = 499)) or
								((vState = 29) and (hState = 500)) or
								((vState = 29) and (hState = 501)) or
								((vState = 29) and (hState = 502)) or
								((vState = 29) and (hState = 510)) or
								((vState = 29) and (hState = 519)) or
								((vState = 29) and (hState = 572)) or
								((vState = 29) and (hState = 576)) or
								((vState = 29) and (hState = 577)) or
								((vState = 29) and (hState = 578)) or
								((vState = 29) and (hState = 579)) or
								((vState = 29) and (hState = 584)) or
								((vState = 29) and (hState = 585)) or
								((vState = 29) and (hState = 586)) or
								((vState = 29) and (hState = 587)) or
								((vState = 29) and (hState = 595)) or
								((vState = 29) and (hState = 596)) or
								((vState = 30) and (hState = 483)) or
								((vState = 30) and (hState = 484)) or
								((vState = 30) and (hState = 485)) or
								((vState = 30) and (hState = 486)) or
								((vState = 30) and (hState = 487)) or
								((vState = 30) and (hState = 488)) or
								((vState = 30) and (hState = 489)) or
								((vState = 30) and (hState = 490)) or
								((vState = 30) and (hState = 491)) or
								((vState = 30) and (hState = 493)) or
								((vState = 30) and (hState = 494)) or
								((vState = 30) and (hState = 495)) or
								((vState = 30) and (hState = 496)) or
								((vState = 30) and (hState = 497)) or
								((vState = 30) and (hState = 498)) or
								((vState = 30) and (hState = 499)) or
								((vState = 30) and (hState = 500)) or
								((vState = 30) and (hState = 501)) or
								((vState = 30) and (hState = 502)) or
								((vState = 30) and (hState = 503)) or
								((vState = 30) and (hState = 510)) or
								((vState = 30) and (hState = 511)) or
								((vState = 30) and (hState = 512)) or
								((vState = 30) and (hState = 518)) or
								((vState = 30) and (hState = 519)) or
								((vState = 30) and (hState = 520)) or
								((vState = 30) and (hState = 572)) or
								((vState = 30) and (hState = 573)) or
								((vState = 30) and (hState = 575)) or
								((vState = 30) and (hState = 576)) or
								((vState = 30) and (hState = 577)) or
								((vState = 30) and (hState = 578)) or
								((vState = 30) and (hState = 579)) or
								((vState = 30) and (hState = 584)) or
								((vState = 30) and (hState = 585)) or
								((vState = 30) and (hState = 586)) or
								((vState = 30) and (hState = 587)) or
								((vState = 30) and (hState = 596)) or
								((vState = 31) and (hState = 482)) or
								((vState = 31) and (hState = 483)) or
								((vState = 31) and (hState = 484)) or
								((vState = 31) and (hState = 485)) or
								((vState = 31) and (hState = 488)) or
								((vState = 31) and (hState = 489)) or
								((vState = 31) and (hState = 490)) or
								((vState = 31) and (hState = 494)) or
								((vState = 31) and (hState = 495)) or
								((vState = 31) and (hState = 496)) or
								((vState = 31) and (hState = 497)) or
								((vState = 31) and (hState = 500)) or
								((vState = 31) and (hState = 501)) or
								((vState = 31) and (hState = 502)) or
								((vState = 31) and (hState = 503)) or
								((vState = 31) and (hState = 504)) or
								((vState = 31) and (hState = 511)) or
								((vState = 31) and (hState = 512)) or
								((vState = 31) and (hState = 513)) or
								((vState = 31) and (hState = 519)) or
								((vState = 31) and (hState = 520)) or
								((vState = 31) and (hState = 572)) or
								((vState = 31) and (hState = 573)) or
								((vState = 31) and (hState = 575)) or
								((vState = 31) and (hState = 576)) or
								((vState = 31) and (hState = 577)) or
								((vState = 31) and (hState = 578)) or
								((vState = 31) and (hState = 579)) or
								((vState = 31) and (hState = 582)) or
								((vState = 31) and (hState = 583)) or
								((vState = 31) and (hState = 584)) or
								((vState = 31) and (hState = 585)) or
								((vState = 31) and (hState = 586)) or
								((vState = 31) and (hState = 587)) or
								((vState = 31) and (hState = 596)) or
								((vState = 31) and (hState = 597)) or
								((vState = 32) and (hState = 480)) or
								((vState = 32) and (hState = 481)) or
								((vState = 32) and (hState = 482)) or
								((vState = 32) and (hState = 483)) or
								((vState = 32) and (hState = 487)) or
								((vState = 32) and (hState = 488)) or
								((vState = 32) and (hState = 489)) or
								((vState = 32) and (hState = 493)) or
								((vState = 32) and (hState = 494)) or
								((vState = 32) and (hState = 495)) or
								((vState = 32) and (hState = 496)) or
								((vState = 32) and (hState = 497)) or
								((vState = 32) and (hState = 498)) or
								((vState = 32) and (hState = 499)) or
								((vState = 32) and (hState = 500)) or
								((vState = 32) and (hState = 503)) or
								((vState = 32) and (hState = 504)) or
								((vState = 32) and (hState = 505)) or
								((vState = 32) and (hState = 506)) or
								((vState = 32) and (hState = 512)) or
								((vState = 32) and (hState = 513)) or
								((vState = 32) and (hState = 514)) or
								((vState = 32) and (hState = 515)) or
								((vState = 32) and (hState = 520)) or
								((vState = 32) and (hState = 521)) or
								((vState = 32) and (hState = 572)) or
								((vState = 32) and (hState = 573)) or
								((vState = 32) and (hState = 575)) or
								((vState = 32) and (hState = 576)) or
								((vState = 32) and (hState = 578)) or
								((vState = 32) and (hState = 579)) or
								((vState = 32) and (hState = 580)) or
								((vState = 32) and (hState = 582)) or
								((vState = 32) and (hState = 583)) or
								((vState = 32) and (hState = 584)) or
								((vState = 32) and (hState = 585)) or
								((vState = 32) and (hState = 586)) or
								((vState = 32) and (hState = 587)) or
								((vState = 32) and (hState = 588)) or
								((vState = 32) and (hState = 589)) or
								((vState = 32) and (hState = 590)) or
								((vState = 32) and (hState = 591)) or
								((vState = 32) and (hState = 592)) or
								((vState = 32) and (hState = 593)) or
								((vState = 32) and (hState = 594)) or
								((vState = 32) and (hState = 596)) or
								((vState = 32) and (hState = 597)) or
								((vState = 33) and (hState = 475)) or
								((vState = 33) and (hState = 476)) or
								((vState = 33) and (hState = 477)) or
								((vState = 33) and (hState = 478)) or
								((vState = 33) and (hState = 479)) or
								((vState = 33) and (hState = 480)) or
								((vState = 33) and (hState = 481)) or
								((vState = 33) and (hState = 482)) or
								((vState = 33) and (hState = 483)) or
								((vState = 33) and (hState = 486)) or
								((vState = 33) and (hState = 487)) or
								((vState = 33) and (hState = 488)) or
								((vState = 33) and (hState = 491)) or
								((vState = 33) and (hState = 492)) or
								((vState = 33) and (hState = 493)) or
								((vState = 33) and (hState = 494)) or
								((vState = 33) and (hState = 497)) or
								((vState = 33) and (hState = 498)) or
								((vState = 33) and (hState = 499)) or
								((vState = 33) and (hState = 500)) or
								((vState = 33) and (hState = 501)) or
								((vState = 33) and (hState = 505)) or
								((vState = 33) and (hState = 506)) or
								((vState = 33) and (hState = 507)) or
								((vState = 33) and (hState = 508)) or
								((vState = 33) and (hState = 509)) or
								((vState = 33) and (hState = 514)) or
								((vState = 33) and (hState = 515)) or
								((vState = 33) and (hState = 516)) or
								((vState = 33) and (hState = 517)) or
								((vState = 33) and (hState = 520)) or
								((vState = 33) and (hState = 521)) or
								((vState = 33) and (hState = 522)) or
								((vState = 33) and (hState = 572)) or
								((vState = 33) and (hState = 573)) or
								((vState = 33) and (hState = 575)) or
								((vState = 33) and (hState = 576)) or
								((vState = 33) and (hState = 579)) or
								((vState = 33) and (hState = 580)) or
								((vState = 33) and (hState = 581)) or
								((vState = 33) and (hState = 582)) or
								((vState = 33) and (hState = 583)) or
								((vState = 33) and (hState = 584)) or
								((vState = 33) and (hState = 585)) or
								((vState = 33) and (hState = 591)) or
								((vState = 33) and (hState = 592)) or
								((vState = 33) and (hState = 593)) or
								((vState = 33) and (hState = 594)) or
								((vState = 33) and (hState = 595)) or
								((vState = 33) and (hState = 596)) or
								((vState = 33) and (hState = 597)) or
								((vState = 34) and (hState = 475)) or
								((vState = 34) and (hState = 476)) or
								((vState = 34) and (hState = 477)) or
								((vState = 34) and (hState = 478)) or
								((vState = 34) and (hState = 479)) or
								((vState = 34) and (hState = 480)) or
								((vState = 34) and (hState = 481)) or
								((vState = 34) and (hState = 482)) or
								((vState = 34) and (hState = 483)) or
								((vState = 34) and (hState = 484)) or
								((vState = 34) and (hState = 485)) or
								((vState = 34) and (hState = 486)) or
								((vState = 34) and (hState = 487)) or
								((vState = 34) and (hState = 488)) or
								((vState = 34) and (hState = 489)) or
								((vState = 34) and (hState = 490)) or
								((vState = 34) and (hState = 491)) or
								((vState = 34) and (hState = 492)) or
								((vState = 34) and (hState = 493)) or
								((vState = 34) and (hState = 497)) or
								((vState = 34) and (hState = 498)) or
								((vState = 34) and (hState = 499)) or
								((vState = 34) and (hState = 500)) or
								((vState = 34) and (hState = 501)) or
								((vState = 34) and (hState = 502)) or
								((vState = 34) and (hState = 503)) or
								((vState = 34) and (hState = 504)) or
								((vState = 34) and (hState = 505)) or
								((vState = 34) and (hState = 506)) or
								((vState = 34) and (hState = 507)) or
								((vState = 34) and (hState = 508)) or
								((vState = 34) and (hState = 509)) or
								((vState = 34) and (hState = 510)) or
								((vState = 34) and (hState = 511)) or
								((vState = 34) and (hState = 512)) or
								((vState = 34) and (hState = 513)) or
								((vState = 34) and (hState = 516)) or
								((vState = 34) and (hState = 517)) or
								((vState = 34) and (hState = 518)) or
								((vState = 34) and (hState = 519)) or
								((vState = 34) and (hState = 521)) or
								((vState = 34) and (hState = 522)) or
								((vState = 34) and (hState = 523)) or
								((vState = 34) and (hState = 570)) or
								((vState = 34) and (hState = 572)) or
								((vState = 34) and (hState = 573)) or
								((vState = 34) and (hState = 574)) or
								((vState = 34) and (hState = 575)) or
								((vState = 34) and (hState = 576)) or
								((vState = 34) and (hState = 580)) or
								((vState = 34) and (hState = 581)) or
								((vState = 34) and (hState = 582)) or
								((vState = 34) and (hState = 583)) or
								((vState = 34) and (hState = 584)) or
								((vState = 34) and (hState = 585)) or
								((vState = 34) and (hState = 590)) or
								((vState = 34) and (hState = 591)) or
								((vState = 34) and (hState = 592)) or
								((vState = 34) and (hState = 593)) or
								((vState = 34) and (hState = 594)) or
								((vState = 34) and (hState = 595)) or
								((vState = 34) and (hState = 596)) or
								((vState = 34) and (hState = 597)) or
								((vState = 34) and (hState = 598)) or
								((vState = 35) and (hState = 475)) or
								((vState = 35) and (hState = 476)) or
								((vState = 35) and (hState = 477)) or
								((vState = 35) and (hState = 478)) or
								((vState = 35) and (hState = 483)) or
								((vState = 35) and (hState = 484)) or
								((vState = 35) and (hState = 485)) or
								((vState = 35) and (hState = 486)) or
								((vState = 35) and (hState = 487)) or
								((vState = 35) and (hState = 488)) or
								((vState = 35) and (hState = 489)) or
								((vState = 35) and (hState = 490)) or
								((vState = 35) and (hState = 491)) or
								((vState = 35) and (hState = 492)) or
								((vState = 35) and (hState = 493)) or
								((vState = 35) and (hState = 497)) or
								((vState = 35) and (hState = 498)) or
								((vState = 35) and (hState = 502)) or
								((vState = 35) and (hState = 503)) or
								((vState = 35) and (hState = 504)) or
								((vState = 35) and (hState = 505)) or
								((vState = 35) and (hState = 506)) or
								((vState = 35) and (hState = 507)) or
								((vState = 35) and (hState = 508)) or
								((vState = 35) and (hState = 509)) or
								((vState = 35) and (hState = 510)) or
								((vState = 35) and (hState = 511)) or
								((vState = 35) and (hState = 512)) or
								((vState = 35) and (hState = 513)) or
								((vState = 35) and (hState = 518)) or
								((vState = 35) and (hState = 519)) or
								((vState = 35) and (hState = 520)) or
								((vState = 35) and (hState = 522)) or
								((vState = 35) and (hState = 523)) or
								((vState = 35) and (hState = 524)) or
								((vState = 35) and (hState = 570)) or
								((vState = 35) and (hState = 571)) or
								((vState = 35) and (hState = 572)) or
								((vState = 35) and (hState = 573)) or
								((vState = 35) and (hState = 574)) or
								((vState = 35) and (hState = 575)) or
								((vState = 35) and (hState = 576)) or
								((vState = 35) and (hState = 581)) or
								((vState = 35) and (hState = 582)) or
								((vState = 35) and (hState = 583)) or
								((vState = 35) and (hState = 584)) or
								((vState = 35) and (hState = 587)) or
								((vState = 35) and (hState = 588)) or
								((vState = 35) and (hState = 589)) or
								((vState = 35) and (hState = 590)) or
								((vState = 35) and (hState = 591)) or
								((vState = 35) and (hState = 592)) or
								((vState = 35) and (hState = 597)) or
								((vState = 35) and (hState = 598)) or
								((vState = 35) and (hState = 599)) or
								((vState = 36) and (hState = 473)) or
								((vState = 36) and (hState = 474)) or
								((vState = 36) and (hState = 475)) or
								((vState = 36) and (hState = 476)) or
								((vState = 36) and (hState = 483)) or
								((vState = 36) and (hState = 484)) or
								((vState = 36) and (hState = 487)) or
								((vState = 36) and (hState = 488)) or
								((vState = 36) and (hState = 489)) or
								((vState = 36) and (hState = 490)) or
								((vState = 36) and (hState = 491)) or
								((vState = 36) and (hState = 492)) or
								((vState = 36) and (hState = 493)) or
								((vState = 36) and (hState = 494)) or
								((vState = 36) and (hState = 495)) or
								((vState = 36) and (hState = 496)) or
								((vState = 36) and (hState = 497)) or
								((vState = 36) and (hState = 498)) or
								((vState = 36) and (hState = 499)) or
								((vState = 36) and (hState = 500)) or
								((vState = 36) and (hState = 501)) or
								((vState = 36) and (hState = 502)) or
								((vState = 36) and (hState = 503)) or
								((vState = 36) and (hState = 504)) or
								((vState = 36) and (hState = 505)) or
								((vState = 36) and (hState = 506)) or
								((vState = 36) and (hState = 507)) or
								((vState = 36) and (hState = 508)) or
								((vState = 36) and (hState = 509)) or
								((vState = 36) and (hState = 510)) or
								((vState = 36) and (hState = 511)) or
								((vState = 36) and (hState = 512)) or
								((vState = 36) and (hState = 513)) or
								((vState = 36) and (hState = 514)) or
								((vState = 36) and (hState = 515)) or
								((vState = 36) and (hState = 516)) or
								((vState = 36) and (hState = 519)) or
								((vState = 36) and (hState = 520)) or
								((vState = 36) and (hState = 521)) or
								((vState = 36) and (hState = 522)) or
								((vState = 36) and (hState = 523)) or
								((vState = 36) and (hState = 524)) or
								((vState = 36) and (hState = 525)) or
								((vState = 36) and (hState = 570)) or
								((vState = 36) and (hState = 571)) or
								((vState = 36) and (hState = 572)) or
								((vState = 36) and (hState = 573)) or
								((vState = 36) and (hState = 574)) or
								((vState = 36) and (hState = 575)) or
								((vState = 36) and (hState = 576)) or
								((vState = 36) and (hState = 582)) or
								((vState = 36) and (hState = 583)) or
								((vState = 36) and (hState = 584)) or
								((vState = 36) and (hState = 585)) or
								((vState = 36) and (hState = 586)) or
								((vState = 36) and (hState = 587)) or
								((vState = 36) and (hState = 588)) or
								((vState = 36) and (hState = 589)) or
								((vState = 36) and (hState = 597)) or
								((vState = 36) and (hState = 598)) or
								((vState = 36) and (hState = 599)) or
								((vState = 37) and (hState = 472)) or
								((vState = 37) and (hState = 473)) or
								((vState = 37) and (hState = 474)) or
								((vState = 37) and (hState = 475)) or
								((vState = 37) and (hState = 476)) or
								((vState = 37) and (hState = 482)) or
								((vState = 37) and (hState = 483)) or
								((vState = 37) and (hState = 486)) or
								((vState = 37) and (hState = 487)) or
								((vState = 37) and (hState = 488)) or
								((vState = 37) and (hState = 489)) or
								((vState = 37) and (hState = 490)) or
								((vState = 37) and (hState = 491)) or
								((vState = 37) and (hState = 494)) or
								((vState = 37) and (hState = 495)) or
								((vState = 37) and (hState = 496)) or
								((vState = 37) and (hState = 497)) or
								((vState = 37) and (hState = 498)) or
								((vState = 37) and (hState = 499)) or
								((vState = 37) and (hState = 500)) or
								((vState = 37) and (hState = 511)) or
								((vState = 37) and (hState = 512)) or
								((vState = 37) and (hState = 513)) or
								((vState = 37) and (hState = 514)) or
								((vState = 37) and (hState = 515)) or
								((vState = 37) and (hState = 516)) or
								((vState = 37) and (hState = 517)) or
								((vState = 37) and (hState = 518)) or
								((vState = 37) and (hState = 520)) or
								((vState = 37) and (hState = 521)) or
								((vState = 37) and (hState = 522)) or
								((vState = 37) and (hState = 523)) or
								((vState = 37) and (hState = 524)) or
								((vState = 37) and (hState = 525)) or
								((vState = 37) and (hState = 526)) or
								((vState = 37) and (hState = 571)) or
								((vState = 37) and (hState = 572)) or
								((vState = 37) and (hState = 573)) or
								((vState = 37) and (hState = 574)) or
								((vState = 37) and (hState = 575)) or
								((vState = 37) and (hState = 576)) or
								((vState = 37) and (hState = 581)) or
								((vState = 37) and (hState = 582)) or
								((vState = 37) and (hState = 583)) or
								((vState = 37) and (hState = 584)) or
								((vState = 37) and (hState = 585)) or
								((vState = 37) and (hState = 586)) or
								((vState = 37) and (hState = 587)) or
								((vState = 37) and (hState = 588)) or
								((vState = 37) and (hState = 589)) or
								((vState = 37) and (hState = 598)) or
								((vState = 38) and (hState = 470)) or
								((vState = 38) and (hState = 471)) or
								((vState = 38) and (hState = 472)) or
								((vState = 38) and (hState = 473)) or
								((vState = 38) and (hState = 475)) or
								((vState = 38) and (hState = 476)) or
								((vState = 38) and (hState = 480)) or
								((vState = 38) and (hState = 481)) or
								((vState = 38) and (hState = 482)) or
								((vState = 38) and (hState = 483)) or
								((vState = 38) and (hState = 484)) or
								((vState = 38) and (hState = 485)) or
								((vState = 38) and (hState = 486)) or
								((vState = 38) and (hState = 487)) or
								((vState = 38) and (hState = 488)) or
								((vState = 38) and (hState = 495)) or
								((vState = 38) and (hState = 496)) or
								((vState = 38) and (hState = 497)) or
								((vState = 38) and (hState = 498)) or
								((vState = 38) and (hState = 499)) or
								((vState = 38) and (hState = 500)) or
								((vState = 38) and (hState = 512)) or
								((vState = 38) and (hState = 513)) or
								((vState = 38) and (hState = 514)) or
								((vState = 38) and (hState = 515)) or
								((vState = 38) and (hState = 516)) or
								((vState = 38) and (hState = 517)) or
								((vState = 38) and (hState = 518)) or
								((vState = 38) and (hState = 519)) or
								((vState = 38) and (hState = 520)) or
								((vState = 38) and (hState = 521)) or
								((vState = 38) and (hState = 522)) or
								((vState = 38) and (hState = 523)) or
								((vState = 38) and (hState = 524)) or
								((vState = 38) and (hState = 525)) or
								((vState = 38) and (hState = 526)) or
								((vState = 38) and (hState = 527)) or
								((vState = 38) and (hState = 571)) or
								((vState = 38) and (hState = 572)) or
								((vState = 38) and (hState = 573)) or
								((vState = 38) and (hState = 574)) or
								((vState = 38) and (hState = 575)) or
								((vState = 38) and (hState = 576)) or
								((vState = 38) and (hState = 577)) or
								((vState = 38) and (hState = 578)) or
								((vState = 38) and (hState = 579)) or
								((vState = 38) and (hState = 580)) or
								((vState = 38) and (hState = 581)) or
								((vState = 38) and (hState = 582)) or
								((vState = 38) and (hState = 583)) or
								((vState = 38) and (hState = 584)) or
								((vState = 38) and (hState = 585)) or
								((vState = 38) and (hState = 586)) or
								((vState = 38) and (hState = 587)) or
								((vState = 38) and (hState = 588)) or
								((vState = 38) and (hState = 589)) or
								((vState = 38) and (hState = 594)) or
								((vState = 38) and (hState = 595)) or
								((vState = 38) and (hState = 596)) or
								((vState = 38) and (hState = 597)) or
								((vState = 38) and (hState = 598)) or
								((vState = 38) and (hState = 599)) or
								((vState = 39) and (hState = 470)) or
								((vState = 39) and (hState = 471)) or
								((vState = 39) and (hState = 475)) or
								((vState = 39) and (hState = 476)) or
								((vState = 39) and (hState = 479)) or
								((vState = 39) and (hState = 480)) or
								((vState = 39) and (hState = 481)) or
								((vState = 39) and (hState = 482)) or
								((vState = 39) and (hState = 483)) or
								((vState = 39) and (hState = 484)) or
								((vState = 39) and (hState = 485)) or
								((vState = 39) and (hState = 493)) or
								((vState = 39) and (hState = 494)) or
								((vState = 39) and (hState = 495)) or
								((vState = 39) and (hState = 496)) or
								((vState = 39) and (hState = 497)) or
								((vState = 39) and (hState = 498)) or
								((vState = 39) and (hState = 499)) or
								((vState = 39) and (hState = 500)) or
								((vState = 39) and (hState = 501)) or
								((vState = 39) and (hState = 511)) or
								((vState = 39) and (hState = 512)) or
								((vState = 39) and (hState = 513)) or
								((vState = 39) and (hState = 514)) or
								((vState = 39) and (hState = 515)) or
								((vState = 39) and (hState = 518)) or
								((vState = 39) and (hState = 519)) or
								((vState = 39) and (hState = 520)) or
								((vState = 39) and (hState = 521)) or
								((vState = 39) and (hState = 522)) or
								((vState = 39) and (hState = 523)) or
								((vState = 39) and (hState = 524)) or
								((vState = 39) and (hState = 525)) or
								((vState = 39) and (hState = 526)) or
								((vState = 39) and (hState = 527)) or
								((vState = 39) and (hState = 528)) or
								((vState = 39) and (hState = 571)) or
								((vState = 39) and (hState = 572)) or
								((vState = 39) and (hState = 573)) or
								((vState = 39) and (hState = 574)) or
								((vState = 39) and (hState = 575)) or
								((vState = 39) and (hState = 576)) or
								((vState = 39) and (hState = 577)) or
								((vState = 39) and (hState = 578)) or
								((vState = 39) and (hState = 579)) or
								((vState = 39) and (hState = 581)) or
								((vState = 39) and (hState = 582)) or
								((vState = 39) and (hState = 583)) or
								((vState = 39) and (hState = 584)) or
								((vState = 39) and (hState = 586)) or
								((vState = 39) and (hState = 587)) or
								((vState = 39) and (hState = 588)) or
								((vState = 39) and (hState = 589)) or
								((vState = 39) and (hState = 590)) or
								((vState = 39) and (hState = 593)) or
								((vState = 39) and (hState = 594)) or
								((vState = 39) and (hState = 595)) or
								((vState = 40) and (hState = 470)) or
								((vState = 40) and (hState = 471)) or
								((vState = 40) and (hState = 475)) or
								((vState = 40) and (hState = 476)) or
								((vState = 40) and (hState = 478)) or
								((vState = 40) and (hState = 479)) or
								((vState = 40) and (hState = 480)) or
								((vState = 40) and (hState = 481)) or
								((vState = 40) and (hState = 482)) or
								((vState = 40) and (hState = 483)) or
								((vState = 40) and (hState = 491)) or
								((vState = 40) and (hState = 492)) or
								((vState = 40) and (hState = 493)) or
								((vState = 40) and (hState = 494)) or
								((vState = 40) and (hState = 495)) or
								((vState = 40) and (hState = 496)) or
								((vState = 40) and (hState = 497)) or
								((vState = 40) and (hState = 498)) or
								((vState = 40) and (hState = 499)) or
								((vState = 40) and (hState = 500)) or
								((vState = 40) and (hState = 501)) or
								((vState = 40) and (hState = 502)) or
								((vState = 40) and (hState = 503)) or
								((vState = 40) and (hState = 504)) or
								((vState = 40) and (hState = 505)) or
								((vState = 40) and (hState = 506)) or
								((vState = 40) and (hState = 507)) or
								((vState = 40) and (hState = 508)) or
								((vState = 40) and (hState = 509)) or
								((vState = 40) and (hState = 510)) or
								((vState = 40) and (hState = 511)) or
								((vState = 40) and (hState = 512)) or
								((vState = 40) and (hState = 513)) or
								((vState = 40) and (hState = 514)) or
								((vState = 40) and (hState = 523)) or
								((vState = 40) and (hState = 524)) or
								((vState = 40) and (hState = 528)) or
								((vState = 40) and (hState = 529)) or
								((vState = 40) and (hState = 572)) or
								((vState = 40) and (hState = 573)) or
								((vState = 40) and (hState = 574)) or
								((vState = 40) and (hState = 575)) or
								((vState = 40) and (hState = 576)) or
								((vState = 40) and (hState = 577)) or
								((vState = 40) and (hState = 578)) or
								((vState = 40) and (hState = 581)) or
								((vState = 40) and (hState = 582)) or
								((vState = 40) and (hState = 583)) or
								((vState = 40) and (hState = 584)) or
								((vState = 40) and (hState = 587)) or
								((vState = 40) and (hState = 588)) or
								((vState = 40) and (hState = 589)) or
								((vState = 40) and (hState = 590)) or
								((vState = 40) and (hState = 594)) or
								((vState = 40) and (hState = 595)) or
								((vState = 41) and (hState = 470)) or
								((vState = 41) and (hState = 471)) or
								((vState = 41) and (hState = 475)) or
								((vState = 41) and (hState = 476)) or
								((vState = 41) and (hState = 477)) or
								((vState = 41) and (hState = 478)) or
								((vState = 41) and (hState = 479)) or
								((vState = 41) and (hState = 481)) or
								((vState = 41) and (hState = 482)) or
								((vState = 41) and (hState = 487)) or
								((vState = 41) and (hState = 488)) or
								((vState = 41) and (hState = 489)) or
								((vState = 41) and (hState = 490)) or
								((vState = 41) and (hState = 491)) or
								((vState = 41) and (hState = 492)) or
								((vState = 41) and (hState = 493)) or
								((vState = 41) and (hState = 494)) or
								((vState = 41) and (hState = 495)) or
								((vState = 41) and (hState = 496)) or
								((vState = 41) and (hState = 497)) or
								((vState = 41) and (hState = 498)) or
								((vState = 41) and (hState = 499)) or
								((vState = 41) and (hState = 500)) or
								((vState = 41) and (hState = 501)) or
								((vState = 41) and (hState = 502)) or
								((vState = 41) and (hState = 503)) or
								((vState = 41) and (hState = 504)) or
								((vState = 41) and (hState = 505)) or
								((vState = 41) and (hState = 506)) or
								((vState = 41) and (hState = 507)) or
								((vState = 41) and (hState = 508)) or
								((vState = 41) and (hState = 509)) or
								((vState = 41) and (hState = 510)) or
								((vState = 41) and (hState = 511)) or
								((vState = 41) and (hState = 512)) or
								((vState = 41) and (hState = 513)) or
								((vState = 41) and (hState = 524)) or
								((vState = 41) and (hState = 525)) or
								((vState = 41) and (hState = 529)) or
								((vState = 41) and (hState = 530)) or
								((vState = 41) and (hState = 572)) or
								((vState = 41) and (hState = 573)) or
								((vState = 41) and (hState = 574)) or
								((vState = 41) and (hState = 576)) or
								((vState = 41) and (hState = 577)) or
								((vState = 41) and (hState = 578)) or
								((vState = 41) and (hState = 579)) or
								((vState = 41) and (hState = 580)) or
								((vState = 41) and (hState = 581)) or
								((vState = 41) and (hState = 582)) or
								((vState = 41) and (hState = 583)) or
								((vState = 41) and (hState = 584)) or
								((vState = 41) and (hState = 585)) or
								((vState = 41) and (hState = 588)) or
								((vState = 41) and (hState = 589)) or
								((vState = 41) and (hState = 590)) or
								((vState = 41) and (hState = 591)) or
								((vState = 41) and (hState = 594)) or
								((vState = 41) and (hState = 595)) or
								((vState = 42) and (hState = 471)) or
								((vState = 42) and (hState = 472)) or
								((vState = 42) and (hState = 475)) or
								((vState = 42) and (hState = 476)) or
								((vState = 42) and (hState = 477)) or
								((vState = 42) and (hState = 478)) or
								((vState = 42) and (hState = 480)) or
								((vState = 42) and (hState = 481)) or
								((vState = 42) and (hState = 485)) or
								((vState = 42) and (hState = 486)) or
								((vState = 42) and (hState = 487)) or
								((vState = 42) and (hState = 488)) or
								((vState = 42) and (hState = 489)) or
								((vState = 42) and (hState = 490)) or
								((vState = 42) and (hState = 498)) or
								((vState = 42) and (hState = 499)) or
								((vState = 42) and (hState = 500)) or
								((vState = 42) and (hState = 501)) or
								((vState = 42) and (hState = 502)) or
								((vState = 42) and (hState = 503)) or
								((vState = 42) and (hState = 504)) or
								((vState = 42) and (hState = 505)) or
								((vState = 42) and (hState = 511)) or
								((vState = 42) and (hState = 512)) or
								((vState = 42) and (hState = 513)) or
								((vState = 42) and (hState = 514)) or
								((vState = 42) and (hState = 525)) or
								((vState = 42) and (hState = 526)) or
								((vState = 42) and (hState = 530)) or
								((vState = 42) and (hState = 531)) or
								((vState = 42) and (hState = 572)) or
								((vState = 42) and (hState = 573)) or
								((vState = 42) and (hState = 574)) or
								((vState = 42) and (hState = 575)) or
								((vState = 42) and (hState = 576)) or
								((vState = 42) and (hState = 577)) or
								((vState = 42) and (hState = 579)) or
								((vState = 42) and (hState = 580)) or
								((vState = 42) and (hState = 581)) or
								((vState = 42) and (hState = 582)) or
								((vState = 42) and (hState = 583)) or
								((vState = 42) and (hState = 584)) or
								((vState = 42) and (hState = 585)) or
								((vState = 42) and (hState = 589)) or
								((vState = 42) and (hState = 590)) or
								((vState = 42) and (hState = 591)) or
								((vState = 42) and (hState = 592)) or
								((vState = 42) and (hState = 594)) or
								((vState = 42) and (hState = 595)) or
								((vState = 43) and (hState = 471)) or
								((vState = 43) and (hState = 472)) or
								((vState = 43) and (hState = 475)) or
								((vState = 43) and (hState = 476)) or
								((vState = 43) and (hState = 477)) or
								((vState = 43) and (hState = 478)) or
								((vState = 43) and (hState = 479)) or
								((vState = 43) and (hState = 480)) or
								((vState = 43) and (hState = 481)) or
								((vState = 43) and (hState = 483)) or
								((vState = 43) and (hState = 484)) or
								((vState = 43) and (hState = 485)) or
								((vState = 43) and (hState = 486)) or
								((vState = 43) and (hState = 487)) or
								((vState = 43) and (hState = 488)) or
								((vState = 43) and (hState = 489)) or
								((vState = 43) and (hState = 498)) or
								((vState = 43) and (hState = 499)) or
								((vState = 43) and (hState = 500)) or
								((vState = 43) and (hState = 501)) or
								((vState = 43) and (hState = 502)) or
								((vState = 43) and (hState = 503)) or
								((vState = 43) and (hState = 504)) or
								((vState = 43) and (hState = 505)) or
								((vState = 43) and (hState = 511)) or
								((vState = 43) and (hState = 512)) or
								((vState = 43) and (hState = 513)) or
								((vState = 43) and (hState = 514)) or
								((vState = 43) and (hState = 515)) or
								((vState = 43) and (hState = 525)) or
								((vState = 43) and (hState = 526)) or
								((vState = 43) and (hState = 527)) or
								((vState = 43) and (hState = 531)) or
								((vState = 43) and (hState = 532)) or
								((vState = 43) and (hState = 572)) or
								((vState = 43) and (hState = 573)) or
								((vState = 43) and (hState = 574)) or
								((vState = 43) and (hState = 575)) or
								((vState = 43) and (hState = 576)) or
								((vState = 43) and (hState = 577)) or
								((vState = 43) and (hState = 580)) or
								((vState = 43) and (hState = 581)) or
								((vState = 43) and (hState = 582)) or
								((vState = 43) and (hState = 583)) or
								((vState = 43) and (hState = 584)) or
								((vState = 43) and (hState = 585)) or
								((vState = 43) and (hState = 589)) or
								((vState = 43) and (hState = 590)) or
								((vState = 43) and (hState = 591)) or
								((vState = 43) and (hState = 592)) or
								((vState = 43) and (hState = 593)) or
								((vState = 43) and (hState = 594)) or
								((vState = 43) and (hState = 595)) or
								((vState = 43) and (hState = 596)) or
								((vState = 44) and (hState = 471)) or
								((vState = 44) and (hState = 472)) or
								((vState = 44) and (hState = 475)) or
								((vState = 44) and (hState = 476)) or
								((vState = 44) and (hState = 477)) or
								((vState = 44) and (hState = 478)) or
								((vState = 44) and (hState = 479)) or
								((vState = 44) and (hState = 480)) or
								((vState = 44) and (hState = 482)) or
								((vState = 44) and (hState = 483)) or
								((vState = 44) and (hState = 484)) or
								((vState = 44) and (hState = 485)) or
								((vState = 44) and (hState = 486)) or
								((vState = 44) and (hState = 487)) or
								((vState = 44) and (hState = 493)) or
								((vState = 44) and (hState = 494)) or
								((vState = 44) and (hState = 495)) or
								((vState = 44) and (hState = 496)) or
								((vState = 44) and (hState = 497)) or
								((vState = 44) and (hState = 498)) or
								((vState = 44) and (hState = 499)) or
								((vState = 44) and (hState = 500)) or
								((vState = 44) and (hState = 503)) or
								((vState = 44) and (hState = 504)) or
								((vState = 44) and (hState = 505)) or
								((vState = 44) and (hState = 506)) or
								((vState = 44) and (hState = 509)) or
								((vState = 44) and (hState = 510)) or
								((vState = 44) and (hState = 511)) or
								((vState = 44) and (hState = 512)) or
								((vState = 44) and (hState = 513)) or
								((vState = 44) and (hState = 514)) or
								((vState = 44) and (hState = 515)) or
								((vState = 44) and (hState = 516)) or
								((vState = 44) and (hState = 517)) or
								((vState = 44) and (hState = 518)) or
								((vState = 44) and (hState = 519)) or
								((vState = 44) and (hState = 520)) or
								((vState = 44) and (hState = 521)) or
								((vState = 44) and (hState = 525)) or
								((vState = 44) and (hState = 526)) or
								((vState = 44) and (hState = 527)) or
								((vState = 44) and (hState = 528)) or
								((vState = 44) and (hState = 532)) or
								((vState = 44) and (hState = 533)) or
								((vState = 44) and (hState = 572)) or
								((vState = 44) and (hState = 573)) or
								((vState = 44) and (hState = 574)) or
								((vState = 44) and (hState = 575)) or
								((vState = 44) and (hState = 577)) or
								((vState = 44) and (hState = 579)) or
								((vState = 44) and (hState = 580)) or
								((vState = 44) and (hState = 581)) or
								((vState = 44) and (hState = 582)) or
								((vState = 44) and (hState = 583)) or
								((vState = 44) and (hState = 584)) or
								((vState = 44) and (hState = 585)) or
								((vState = 44) and (hState = 589)) or
								((vState = 44) and (hState = 590)) or
								((vState = 44) and (hState = 591)) or
								((vState = 44) and (hState = 592)) or
								((vState = 44) and (hState = 593)) or
								((vState = 44) and (hState = 594)) or
								((vState = 44) and (hState = 595)) or
								((vState = 44) and (hState = 596)) or
								((vState = 45) and (hState = 471)) or
								((vState = 45) and (hState = 472)) or
								((vState = 45) and (hState = 475)) or
								((vState = 45) and (hState = 476)) or
								((vState = 45) and (hState = 477)) or
								((vState = 45) and (hState = 478)) or
								((vState = 45) and (hState = 479)) or
								((vState = 45) and (hState = 480)) or
								((vState = 45) and (hState = 481)) or
								((vState = 45) and (hState = 482)) or
								((vState = 45) and (hState = 483)) or
								((vState = 45) and (hState = 484)) or
								((vState = 45) and (hState = 486)) or
								((vState = 45) and (hState = 487)) or
								((vState = 45) and (hState = 492)) or
								((vState = 45) and (hState = 493)) or
								((vState = 45) and (hState = 494)) or
								((vState = 45) and (hState = 495)) or
								((vState = 45) and (hState = 496)) or
								((vState = 45) and (hState = 497)) or
								((vState = 45) and (hState = 498)) or
								((vState = 45) and (hState = 499)) or
								((vState = 45) and (hState = 500)) or
								((vState = 45) and (hState = 501)) or
								((vState = 45) and (hState = 502)) or
								((vState = 45) and (hState = 503)) or
								((vState = 45) and (hState = 504)) or
								((vState = 45) and (hState = 505)) or
								((vState = 45) and (hState = 506)) or
								((vState = 45) and (hState = 507)) or
								((vState = 45) and (hState = 508)) or
								((vState = 45) and (hState = 509)) or
								((vState = 45) and (hState = 510)) or
								((vState = 45) and (hState = 511)) or
								((vState = 45) and (hState = 512)) or
								((vState = 45) and (hState = 513)) or
								((vState = 45) and (hState = 514)) or
								((vState = 45) and (hState = 515)) or
								((vState = 45) and (hState = 516)) or
								((vState = 45) and (hState = 517)) or
								((vState = 45) and (hState = 518)) or
								((vState = 45) and (hState = 519)) or
								((vState = 45) and (hState = 520)) or
								((vState = 45) and (hState = 521)) or
								((vState = 45) and (hState = 522)) or
								((vState = 45) and (hState = 524)) or
								((vState = 45) and (hState = 525)) or
								((vState = 45) and (hState = 527)) or
								((vState = 45) and (hState = 528)) or
								((vState = 45) and (hState = 529)) or
								((vState = 45) and (hState = 533)) or
								((vState = 45) and (hState = 534)) or
								((vState = 45) and (hState = 573)) or
								((vState = 45) and (hState = 574)) or
								((vState = 45) and (hState = 575)) or
								((vState = 45) and (hState = 576)) or
								((vState = 45) and (hState = 577)) or
								((vState = 45) and (hState = 578)) or
								((vState = 45) and (hState = 579)) or
								((vState = 45) and (hState = 580)) or
								((vState = 45) and (hState = 583)) or
								((vState = 45) and (hState = 584)) or
								((vState = 45) and (hState = 585)) or
								((vState = 45) and (hState = 589)) or
								((vState = 45) and (hState = 590)) or
								((vState = 45) and (hState = 592)) or
								((vState = 45) and (hState = 593)) or
								((vState = 45) and (hState = 594)) or
								((vState = 45) and (hState = 595)) or
								((vState = 45) and (hState = 596)) or
								((vState = 46) and (hState = 472)) or
								((vState = 46) and (hState = 473)) or
								((vState = 46) and (hState = 475)) or
								((vState = 46) and (hState = 476)) or
								((vState = 46) and (hState = 477)) or
								((vState = 46) and (hState = 478)) or
								((vState = 46) and (hState = 479)) or
								((vState = 46) and (hState = 480)) or
								((vState = 46) and (hState = 481)) or
								((vState = 46) and (hState = 482)) or
								((vState = 46) and (hState = 483)) or
								((vState = 46) and (hState = 486)) or
								((vState = 46) and (hState = 487)) or
								((vState = 46) and (hState = 491)) or
								((vState = 46) and (hState = 492)) or
								((vState = 46) and (hState = 493)) or
								((vState = 46) and (hState = 494)) or
								((vState = 46) and (hState = 495)) or
								((vState = 46) and (hState = 496)) or
								((vState = 46) and (hState = 497)) or
								((vState = 46) and (hState = 498)) or
								((vState = 46) and (hState = 500)) or
								((vState = 46) and (hState = 501)) or
								((vState = 46) and (hState = 502)) or
								((vState = 46) and (hState = 503)) or
								((vState = 46) and (hState = 504)) or
								((vState = 46) and (hState = 505)) or
								((vState = 46) and (hState = 506)) or
								((vState = 46) and (hState = 507)) or
								((vState = 46) and (hState = 508)) or
								((vState = 46) and (hState = 509)) or
								((vState = 46) and (hState = 510)) or
								((vState = 46) and (hState = 511)) or
								((vState = 46) and (hState = 512)) or
								((vState = 46) and (hState = 513)) or
								((vState = 46) and (hState = 518)) or
								((vState = 46) and (hState = 519)) or
								((vState = 46) and (hState = 520)) or
								((vState = 46) and (hState = 521)) or
								((vState = 46) and (hState = 522)) or
								((vState = 46) and (hState = 523)) or
								((vState = 46) and (hState = 524)) or
								((vState = 46) and (hState = 525)) or
								((vState = 46) and (hState = 528)) or
								((vState = 46) and (hState = 529)) or
								((vState = 46) and (hState = 530)) or
								((vState = 46) and (hState = 534)) or
								((vState = 46) and (hState = 535)) or
								((vState = 46) and (hState = 568)) or
								((vState = 46) and (hState = 569)) or
								((vState = 46) and (hState = 570)) or
								((vState = 46) and (hState = 571)) or
								((vState = 46) and (hState = 572)) or
								((vState = 46) and (hState = 573)) or
								((vState = 46) and (hState = 574)) or
								((vState = 46) and (hState = 575)) or
								((vState = 46) and (hState = 576)) or
								((vState = 46) and (hState = 577)) or
								((vState = 46) and (hState = 578)) or
								((vState = 46) and (hState = 579)) or
								((vState = 46) and (hState = 584)) or
								((vState = 46) and (hState = 585)) or
								((vState = 46) and (hState = 586)) or
								((vState = 46) and (hState = 587)) or
								((vState = 46) and (hState = 590)) or
								((vState = 46) and (hState = 593)) or
								((vState = 46) and (hState = 594)) or
								((vState = 46) and (hState = 595)) or
								((vState = 46) and (hState = 596)) or
								((vState = 46) and (hState = 597)) or
								((vState = 47) and (hState = 472)) or
								((vState = 47) and (hState = 473)) or
								((vState = 47) and (hState = 475)) or
								((vState = 47) and (hState = 476)) or
								((vState = 47) and (hState = 477)) or
								((vState = 47) and (hState = 478)) or
								((vState = 47) and (hState = 479)) or
								((vState = 47) and (hState = 481)) or
								((vState = 47) and (hState = 482)) or
								((vState = 47) and (hState = 483)) or
								((vState = 47) and (hState = 486)) or
								((vState = 47) and (hState = 487)) or
								((vState = 47) and (hState = 490)) or
								((vState = 47) and (hState = 491)) or
								((vState = 47) and (hState = 492)) or
								((vState = 47) and (hState = 493)) or
								((vState = 47) and (hState = 496)) or
								((vState = 47) and (hState = 497)) or
								((vState = 47) and (hState = 503)) or
								((vState = 47) and (hState = 504)) or
								((vState = 47) and (hState = 505)) or
								((vState = 47) and (hState = 506)) or
								((vState = 47) and (hState = 507)) or
								((vState = 47) and (hState = 508)) or
								((vState = 47) and (hState = 509)) or
								((vState = 47) and (hState = 510)) or
								((vState = 47) and (hState = 511)) or
								((vState = 47) and (hState = 512)) or
								((vState = 47) and (hState = 520)) or
								((vState = 47) and (hState = 521)) or
								((vState = 47) and (hState = 522)) or
								((vState = 47) and (hState = 523)) or
								((vState = 47) and (hState = 524)) or
								((vState = 47) and (hState = 525)) or
								((vState = 47) and (hState = 526)) or
								((vState = 47) and (hState = 529)) or
								((vState = 47) and (hState = 530)) or
								((vState = 47) and (hState = 535)) or
								((vState = 47) and (hState = 536)) or
								((vState = 47) and (hState = 567)) or
								((vState = 47) and (hState = 568)) or
								((vState = 47) and (hState = 569)) or
								((vState = 47) and (hState = 570)) or
								((vState = 47) and (hState = 571)) or
								((vState = 47) and (hState = 572)) or
								((vState = 47) and (hState = 573)) or
								((vState = 47) and (hState = 574)) or
								((vState = 47) and (hState = 575)) or
								((vState = 47) and (hState = 576)) or
								((vState = 47) and (hState = 577)) or
								((vState = 47) and (hState = 578)) or
								((vState = 47) and (hState = 579)) or
								((vState = 47) and (hState = 584)) or
								((vState = 47) and (hState = 585)) or
								((vState = 47) and (hState = 586)) or
								((vState = 47) and (hState = 587)) or
								((vState = 47) and (hState = 588)) or
								((vState = 47) and (hState = 590)) or
								((vState = 47) and (hState = 591)) or
								((vState = 47) and (hState = 594)) or
								((vState = 47) and (hState = 595)) or
								((vState = 47) and (hState = 596)) or
								((vState = 47) and (hState = 597)) or
								((vState = 47) and (hState = 598)) or
								((vState = 48) and (hState = 472)) or
								((vState = 48) and (hState = 473)) or
								((vState = 48) and (hState = 475)) or
								((vState = 48) and (hState = 476)) or
								((vState = 48) and (hState = 477)) or
								((vState = 48) and (hState = 482)) or
								((vState = 48) and (hState = 486)) or
								((vState = 48) and (hState = 487)) or
								((vState = 48) and (hState = 488)) or
								((vState = 48) and (hState = 489)) or
								((vState = 48) and (hState = 490)) or
								((vState = 48) and (hState = 491)) or
								((vState = 48) and (hState = 495)) or
								((vState = 48) and (hState = 496)) or
								((vState = 48) and (hState = 504)) or
								((vState = 48) and (hState = 505)) or
								((vState = 48) and (hState = 506)) or
								((vState = 48) and (hState = 507)) or
								((vState = 48) and (hState = 508)) or
								((vState = 48) and (hState = 509)) or
								((vState = 48) and (hState = 510)) or
								((vState = 48) and (hState = 511)) or
								((vState = 48) and (hState = 512)) or
								((vState = 48) and (hState = 513)) or
								((vState = 48) and (hState = 514)) or
								((vState = 48) and (hState = 515)) or
								((vState = 48) and (hState = 516)) or
								((vState = 48) and (hState = 517)) or
								((vState = 48) and (hState = 518)) or
								((vState = 48) and (hState = 519)) or
								((vState = 48) and (hState = 520)) or
								((vState = 48) and (hState = 521)) or
								((vState = 48) and (hState = 522)) or
								((vState = 48) and (hState = 523)) or
								((vState = 48) and (hState = 524)) or
								((vState = 48) and (hState = 525)) or
								((vState = 48) and (hState = 526)) or
								((vState = 48) and (hState = 529)) or
								((vState = 48) and (hState = 530)) or
								((vState = 48) and (hState = 535)) or
								((vState = 48) and (hState = 536)) or
								((vState = 48) and (hState = 537)) or
								((vState = 48) and (hState = 565)) or
								((vState = 48) and (hState = 566)) or
								((vState = 48) and (hState = 567)) or
								((vState = 48) and (hState = 568)) or
								((vState = 48) and (hState = 571)) or
								((vState = 48) and (hState = 572)) or
								((vState = 48) and (hState = 573)) or
								((vState = 48) and (hState = 574)) or
								((vState = 48) and (hState = 575)) or
								((vState = 48) and (hState = 576)) or
								((vState = 48) and (hState = 577)) or
								((vState = 48) and (hState = 578)) or
								((vState = 48) and (hState = 579)) or
								((vState = 48) and (hState = 582)) or
								((vState = 48) and (hState = 583)) or
								((vState = 48) and (hState = 584)) or
								((vState = 48) and (hState = 585)) or
								((vState = 48) and (hState = 586)) or
								((vState = 48) and (hState = 587)) or
								((vState = 48) and (hState = 588)) or
								((vState = 48) and (hState = 589)) or
								((vState = 48) and (hState = 590)) or
								((vState = 48) and (hState = 591)) or
								((vState = 48) and (hState = 593)) or
								((vState = 48) and (hState = 594)) or
								((vState = 48) and (hState = 596)) or
								((vState = 48) and (hState = 597)) or
								((vState = 48) and (hState = 598)) or
								((vState = 48) and (hState = 599)) or
								((vState = 49) and (hState = 472)) or
								((vState = 49) and (hState = 473)) or
								((vState = 49) and (hState = 474)) or
								((vState = 49) and (hState = 475)) or
								((vState = 49) and (hState = 476)) or
								((vState = 49) and (hState = 482)) or
								((vState = 49) and (hState = 486)) or
								((vState = 49) and (hState = 487)) or
								((vState = 49) and (hState = 488)) or
								((vState = 49) and (hState = 489)) or
								((vState = 49) and (hState = 490)) or
								((vState = 49) and (hState = 495)) or
								((vState = 49) and (hState = 496)) or
								((vState = 49) and (hState = 498)) or
								((vState = 49) and (hState = 499)) or
								((vState = 49) and (hState = 500)) or
								((vState = 49) and (hState = 501)) or
								((vState = 49) and (hState = 502)) or
								((vState = 49) and (hState = 503)) or
								((vState = 49) and (hState = 504)) or
								((vState = 49) and (hState = 505)) or
								((vState = 49) and (hState = 506)) or
								((vState = 49) and (hState = 508)) or
								((vState = 49) and (hState = 509)) or
								((vState = 49) and (hState = 510)) or
								((vState = 49) and (hState = 511)) or
								((vState = 49) and (hState = 512)) or
								((vState = 49) and (hState = 515)) or
								((vState = 49) and (hState = 516)) or
								((vState = 49) and (hState = 517)) or
								((vState = 49) and (hState = 518)) or
								((vState = 49) and (hState = 519)) or
								((vState = 49) and (hState = 520)) or
								((vState = 49) and (hState = 521)) or
								((vState = 49) and (hState = 522)) or
								((vState = 49) and (hState = 523)) or
								((vState = 49) and (hState = 524)) or
								((vState = 49) and (hState = 525)) or
								((vState = 49) and (hState = 526)) or
								((vState = 49) and (hState = 527)) or
								((vState = 49) and (hState = 529)) or
								((vState = 49) and (hState = 530)) or
								((vState = 49) and (hState = 533)) or
								((vState = 49) and (hState = 534)) or
								((vState = 49) and (hState = 535)) or
								((vState = 49) and (hState = 536)) or
								((vState = 49) and (hState = 537)) or
								((vState = 49) and (hState = 538)) or
								((vState = 49) and (hState = 564)) or
								((vState = 49) and (hState = 565)) or
								((vState = 49) and (hState = 566)) or
								((vState = 49) and (hState = 570)) or
								((vState = 49) and (hState = 571)) or
								((vState = 49) and (hState = 574)) or
								((vState = 49) and (hState = 575)) or
								((vState = 49) and (hState = 576)) or
								((vState = 49) and (hState = 577)) or
								((vState = 49) and (hState = 578)) or
								((vState = 49) and (hState = 579)) or
								((vState = 49) and (hState = 580)) or
								((vState = 49) and (hState = 581)) or
								((vState = 49) and (hState = 582)) or
								((vState = 49) and (hState = 583)) or
								((vState = 49) and (hState = 584)) or
								((vState = 49) and (hState = 585)) or
								((vState = 49) and (hState = 586)) or
								((vState = 49) and (hState = 587)) or
								((vState = 49) and (hState = 588)) or
								((vState = 49) and (hState = 589)) or
								((vState = 49) and (hState = 590)) or
								((vState = 49) and (hState = 591)) or
								((vState = 49) and (hState = 593)) or
								((vState = 49) and (hState = 594)) or
								((vState = 49) and (hState = 598)) or
								((vState = 49) and (hState = 599)) or
								((vState = 50) and (hState = 473)) or
								((vState = 50) and (hState = 474)) or
								((vState = 50) and (hState = 475)) or
								((vState = 50) and (hState = 476)) or
								((vState = 50) and (hState = 482)) or
								((vState = 50) and (hState = 485)) or
								((vState = 50) and (hState = 486)) or
								((vState = 50) and (hState = 487)) or
								((vState = 50) and (hState = 488)) or
								((vState = 50) and (hState = 489)) or
								((vState = 50) and (hState = 490)) or
								((vState = 50) and (hState = 494)) or
								((vState = 50) and (hState = 495)) or
								((vState = 50) and (hState = 496)) or
								((vState = 50) and (hState = 497)) or
								((vState = 50) and (hState = 498)) or
								((vState = 50) and (hState = 499)) or
								((vState = 50) and (hState = 500)) or
								((vState = 50) and (hState = 501)) or
								((vState = 50) and (hState = 502)) or
								((vState = 50) and (hState = 503)) or
								((vState = 50) and (hState = 504)) or
								((vState = 50) and (hState = 505)) or
								((vState = 50) and (hState = 506)) or
								((vState = 50) and (hState = 507)) or
								((vState = 50) and (hState = 508)) or
								((vState = 50) and (hState = 509)) or
								((vState = 50) and (hState = 510)) or
								((vState = 50) and (hState = 511)) or
								((vState = 50) and (hState = 512)) or
								((vState = 50) and (hState = 515)) or
								((vState = 50) and (hState = 516)) or
								((vState = 50) and (hState = 517)) or
								((vState = 50) and (hState = 518)) or
								((vState = 50) and (hState = 519)) or
								((vState = 50) and (hState = 520)) or
								((vState = 50) and (hState = 522)) or
								((vState = 50) and (hState = 523)) or
								((vState = 50) and (hState = 524)) or
								((vState = 50) and (hState = 525)) or
								((vState = 50) and (hState = 526)) or
								((vState = 50) and (hState = 527)) or
								((vState = 50) and (hState = 528)) or
								((vState = 50) and (hState = 529)) or
								((vState = 50) and (hState = 532)) or
								((vState = 50) and (hState = 533)) or
								((vState = 50) and (hState = 534)) or
								((vState = 50) and (hState = 535)) or
								((vState = 50) and (hState = 536)) or
								((vState = 50) and (hState = 537)) or
								((vState = 50) and (hState = 538)) or
								((vState = 50) and (hState = 539)) or
								((vState = 50) and (hState = 562)) or
								((vState = 50) and (hState = 563)) or
								((vState = 50) and (hState = 564)) or
								((vState = 50) and (hState = 569)) or
								((vState = 50) and (hState = 570)) or
								((vState = 50) and (hState = 571)) or
								((vState = 50) and (hState = 574)) or
								((vState = 50) and (hState = 575)) or
								((vState = 50) and (hState = 576)) or
								((vState = 50) and (hState = 577)) or
								((vState = 50) and (hState = 578)) or
								((vState = 50) and (hState = 579)) or
								((vState = 50) and (hState = 580)) or
								((vState = 50) and (hState = 581)) or
								((vState = 50) and (hState = 582)) or
								((vState = 50) and (hState = 583)) or
								((vState = 50) and (hState = 584)) or
								((vState = 50) and (hState = 585)) or
								((vState = 50) and (hState = 586)) or
								((vState = 50) and (hState = 587)) or
								((vState = 50) and (hState = 590)) or
								((vState = 50) and (hState = 591)) or
								((vState = 50) and (hState = 592)) or
								((vState = 50) and (hState = 593)) or
								((vState = 50) and (hState = 594)) or
								((vState = 51) and (hState = 473)) or
								((vState = 51) and (hState = 474)) or
								((vState = 51) and (hState = 475)) or
								((vState = 51) and (hState = 476)) or
								((vState = 51) and (hState = 482)) or
								((vState = 51) and (hState = 484)) or
								((vState = 51) and (hState = 485)) or
								((vState = 51) and (hState = 486)) or
								((vState = 51) and (hState = 487)) or
								((vState = 51) and (hState = 488)) or
								((vState = 51) and (hState = 489)) or
								((vState = 51) and (hState = 494)) or
								((vState = 51) and (hState = 495)) or
								((vState = 51) and (hState = 496)) or
								((vState = 51) and (hState = 497)) or
								((vState = 51) and (hState = 498)) or
								((vState = 51) and (hState = 499)) or
								((vState = 51) and (hState = 500)) or
								((vState = 51) and (hState = 501)) or
								((vState = 51) and (hState = 504)) or
								((vState = 51) and (hState = 505)) or
								((vState = 51) and (hState = 506)) or
								((vState = 51) and (hState = 507)) or
								((vState = 51) and (hState = 508)) or
								((vState = 51) and (hState = 509)) or
								((vState = 51) and (hState = 510)) or
								((vState = 51) and (hState = 511)) or
								((vState = 51) and (hState = 512)) or
								((vState = 51) and (hState = 515)) or
								((vState = 51) and (hState = 516)) or
								((vState = 51) and (hState = 519)) or
								((vState = 51) and (hState = 520)) or
								((vState = 51) and (hState = 521)) or
								((vState = 51) and (hState = 522)) or
								((vState = 51) and (hState = 523)) or
								((vState = 51) and (hState = 525)) or
								((vState = 51) and (hState = 526)) or
								((vState = 51) and (hState = 527)) or
								((vState = 51) and (hState = 528)) or
								((vState = 51) and (hState = 529)) or
								((vState = 51) and (hState = 530)) or
								((vState = 51) and (hState = 531)) or
								((vState = 51) and (hState = 532)) or
								((vState = 51) and (hState = 533)) or
								((vState = 51) and (hState = 536)) or
								((vState = 51) and (hState = 537)) or
								((vState = 51) and (hState = 538)) or
								((vState = 51) and (hState = 539)) or
								((vState = 51) and (hState = 540)) or
								((vState = 51) and (hState = 560)) or
								((vState = 51) and (hState = 561)) or
								((vState = 51) and (hState = 562)) or
								((vState = 51) and (hState = 563)) or
								((vState = 51) and (hState = 568)) or
								((vState = 51) and (hState = 569)) or
								((vState = 51) and (hState = 570)) or
								((vState = 51) and (hState = 571)) or
								((vState = 51) and (hState = 572)) or
								((vState = 51) and (hState = 573)) or
								((vState = 51) and (hState = 574)) or
								((vState = 51) and (hState = 575)) or
								((vState = 51) and (hState = 576)) or
								((vState = 51) and (hState = 577)) or
								((vState = 51) and (hState = 579)) or
								((vState = 51) and (hState = 580)) or
								((vState = 51) and (hState = 584)) or
								((vState = 51) and (hState = 585)) or
								((vState = 51) and (hState = 586)) or
								((vState = 51) and (hState = 587)) or
								((vState = 51) and (hState = 588)) or
								((vState = 51) and (hState = 589)) or
								((vState = 51) and (hState = 590)) or
								((vState = 51) and (hState = 591)) or
								((vState = 51) and (hState = 592)) or
								((vState = 51) and (hState = 593)) or
								((vState = 51) and (hState = 594)) or
								((vState = 52) and (hState = 474)) or
								((vState = 52) and (hState = 475)) or
								((vState = 52) and (hState = 476)) or
								((vState = 52) and (hState = 482)) or
								((vState = 52) and (hState = 484)) or
								((vState = 52) and (hState = 485)) or
								((vState = 52) and (hState = 486)) or
								((vState = 52) and (hState = 487)) or
								((vState = 52) and (hState = 488)) or
								((vState = 52) and (hState = 489)) or
								((vState = 52) and (hState = 493)) or
								((vState = 52) and (hState = 494)) or
								((vState = 52) and (hState = 495)) or
								((vState = 52) and (hState = 496)) or
								((vState = 52) and (hState = 497)) or
								((vState = 52) and (hState = 498)) or
								((vState = 52) and (hState = 499)) or
								((vState = 52) and (hState = 503)) or
								((vState = 52) and (hState = 504)) or
								((vState = 52) and (hState = 505)) or
								((vState = 52) and (hState = 506)) or
								((vState = 52) and (hState = 507)) or
								((vState = 52) and (hState = 508)) or
								((vState = 52) and (hState = 509)) or
								((vState = 52) and (hState = 510)) or
								((vState = 52) and (hState = 511)) or
								((vState = 52) and (hState = 512)) or
								((vState = 52) and (hState = 513)) or
								((vState = 52) and (hState = 514)) or
								((vState = 52) and (hState = 515)) or
								((vState = 52) and (hState = 516)) or
								((vState = 52) and (hState = 521)) or
								((vState = 52) and (hState = 522)) or
								((vState = 52) and (hState = 523)) or
								((vState = 52) and (hState = 526)) or
								((vState = 52) and (hState = 527)) or
								((vState = 52) and (hState = 528)) or
								((vState = 52) and (hState = 529)) or
								((vState = 52) and (hState = 530)) or
								((vState = 52) and (hState = 531)) or
								((vState = 52) and (hState = 532)) or
								((vState = 52) and (hState = 538)) or
								((vState = 52) and (hState = 539)) or
								((vState = 52) and (hState = 540)) or
								((vState = 52) and (hState = 541)) or
								((vState = 52) and (hState = 559)) or
								((vState = 52) and (hState = 560)) or
								((vState = 52) and (hState = 561)) or
								((vState = 52) and (hState = 567)) or
								((vState = 52) and (hState = 568)) or
								((vState = 52) and (hState = 569)) or
								((vState = 52) and (hState = 570)) or
								((vState = 52) and (hState = 571)) or
								((vState = 52) and (hState = 572)) or
								((vState = 52) and (hState = 573)) or
								((vState = 52) and (hState = 574)) or
								((vState = 52) and (hState = 575)) or
								((vState = 52) and (hState = 576)) or
								((vState = 52) and (hState = 577)) or
								((vState = 52) and (hState = 578)) or
								((vState = 52) and (hState = 579)) or
								((vState = 52) and (hState = 580)) or
								((vState = 52) and (hState = 586)) or
								((vState = 52) and (hState = 587)) or
								((vState = 52) and (hState = 588)) or
								((vState = 52) and (hState = 589)) or
								((vState = 52) and (hState = 590)) or
								((vState = 52) and (hState = 591)) or
								((vState = 52) and (hState = 592)) or
								((vState = 52) and (hState = 593)) or
								((vState = 52) and (hState = 594)) or
								((vState = 52) and (hState = 595)) or
								((vState = 53) and (hState = 474)) or
								((vState = 53) and (hState = 475)) or
								((vState = 53) and (hState = 476)) or
								((vState = 53) and (hState = 481)) or
								((vState = 53) and (hState = 482)) or
								((vState = 53) and (hState = 484)) or
								((vState = 53) and (hState = 485)) or
								((vState = 53) and (hState = 486)) or
								((vState = 53) and (hState = 487)) or
								((vState = 53) and (hState = 488)) or
								((vState = 53) and (hState = 489)) or
								((vState = 53) and (hState = 493)) or
								((vState = 53) and (hState = 494)) or
								((vState = 53) and (hState = 495)) or
								((vState = 53) and (hState = 496)) or
								((vState = 53) and (hState = 497)) or
								((vState = 53) and (hState = 503)) or
								((vState = 53) and (hState = 504)) or
								((vState = 53) and (hState = 505)) or
								((vState = 53) and (hState = 506)) or
								((vState = 53) and (hState = 507)) or
								((vState = 53) and (hState = 508)) or
								((vState = 53) and (hState = 509)) or
								((vState = 53) and (hState = 510)) or
								((vState = 53) and (hState = 511)) or
								((vState = 53) and (hState = 512)) or
								((vState = 53) and (hState = 513)) or
								((vState = 53) and (hState = 514)) or
								((vState = 53) and (hState = 515)) or
								((vState = 53) and (hState = 516)) or
								((vState = 53) and (hState = 517)) or
								((vState = 53) and (hState = 518)) or
								((vState = 53) and (hState = 519)) or
								((vState = 53) and (hState = 520)) or
								((vState = 53) and (hState = 521)) or
								((vState = 53) and (hState = 522)) or
								((vState = 53) and (hState = 523)) or
								((vState = 53) and (hState = 524)) or
								((vState = 53) and (hState = 525)) or
								((vState = 53) and (hState = 526)) or
								((vState = 53) and (hState = 527)) or
								((vState = 53) and (hState = 528)) or
								((vState = 53) and (hState = 529)) or
								((vState = 53) and (hState = 530)) or
								((vState = 53) and (hState = 531)) or
								((vState = 53) and (hState = 532)) or
								((vState = 53) and (hState = 533)) or
								((vState = 53) and (hState = 534)) or
								((vState = 53) and (hState = 538)) or
								((vState = 53) and (hState = 539)) or
								((vState = 53) and (hState = 540)) or
								((vState = 53) and (hState = 541)) or
								((vState = 53) and (hState = 542)) or
								((vState = 53) and (hState = 557)) or
								((vState = 53) and (hState = 558)) or
								((vState = 53) and (hState = 559)) or
								((vState = 53) and (hState = 560)) or
								((vState = 53) and (hState = 564)) or
								((vState = 53) and (hState = 565)) or
								((vState = 53) and (hState = 566)) or
								((vState = 53) and (hState = 567)) or
								((vState = 53) and (hState = 568)) or
								((vState = 53) and (hState = 569)) or
								((vState = 53) and (hState = 570)) or
								((vState = 53) and (hState = 571)) or
								((vState = 53) and (hState = 572)) or
								((vState = 53) and (hState = 573)) or
								((vState = 53) and (hState = 574)) or
								((vState = 53) and (hState = 575)) or
								((vState = 53) and (hState = 576)) or
								((vState = 53) and (hState = 577)) or
								((vState = 53) and (hState = 578)) or
								((vState = 53) and (hState = 579)) or
								((vState = 53) and (hState = 580)) or
								((vState = 53) and (hState = 581)) or
								((vState = 53) and (hState = 586)) or
								((vState = 53) and (hState = 587)) or
								((vState = 53) and (hState = 590)) or
								((vState = 53) and (hState = 591)) or
								((vState = 53) and (hState = 592)) or
								((vState = 53) and (hState = 594)) or
								((vState = 53) and (hState = 595)) or
								((vState = 53) and (hState = 596)) or
								((vState = 54) and (hState = 474)) or
								((vState = 54) and (hState = 475)) or
								((vState = 54) and (hState = 481)) or
								((vState = 54) and (hState = 482)) or
								((vState = 54) and (hState = 484)) or
								((vState = 54) and (hState = 485)) or
								((vState = 54) and (hState = 486)) or
								((vState = 54) and (hState = 487)) or
								((vState = 54) and (hState = 488)) or
								((vState = 54) and (hState = 492)) or
								((vState = 54) and (hState = 493)) or
								((vState = 54) and (hState = 494)) or
								((vState = 54) and (hState = 495)) or
								((vState = 54) and (hState = 502)) or
								((vState = 54) and (hState = 503)) or
								((vState = 54) and (hState = 504)) or
								((vState = 54) and (hState = 505)) or
								((vState = 54) and (hState = 506)) or
								((vState = 54) and (hState = 507)) or
								((vState = 54) and (hState = 508)) or
								((vState = 54) and (hState = 509)) or
								((vState = 54) and (hState = 510)) or
								((vState = 54) and (hState = 511)) or
								((vState = 54) and (hState = 512)) or
								((vState = 54) and (hState = 513)) or
								((vState = 54) and (hState = 514)) or
								((vState = 54) and (hState = 515)) or
								((vState = 54) and (hState = 516)) or
								((vState = 54) and (hState = 517)) or
								((vState = 54) and (hState = 518)) or
								((vState = 54) and (hState = 519)) or
								((vState = 54) and (hState = 520)) or
								((vState = 54) and (hState = 521)) or
								((vState = 54) and (hState = 522)) or
								((vState = 54) and (hState = 523)) or
								((vState = 54) and (hState = 524)) or
								((vState = 54) and (hState = 525)) or
								((vState = 54) and (hState = 526)) or
								((vState = 54) and (hState = 527)) or
								((vState = 54) and (hState = 528)) or
								((vState = 54) and (hState = 529)) or
								((vState = 54) and (hState = 533)) or
								((vState = 54) and (hState = 534)) or
								((vState = 54) and (hState = 539)) or
								((vState = 54) and (hState = 540)) or
								((vState = 54) and (hState = 541)) or
								((vState = 54) and (hState = 542)) or
								((vState = 54) and (hState = 543)) or
								((vState = 54) and (hState = 555)) or
								((vState = 54) and (hState = 556)) or
								((vState = 54) and (hState = 557)) or
								((vState = 54) and (hState = 558)) or
								((vState = 54) and (hState = 562)) or
								((vState = 54) and (hState = 563)) or
								((vState = 54) and (hState = 564)) or
								((vState = 54) and (hState = 565)) or
								((vState = 54) and (hState = 566)) or
								((vState = 54) and (hState = 567)) or
								((vState = 54) and (hState = 568)) or
								((vState = 54) and (hState = 569)) or
								((vState = 54) and (hState = 570)) or
								((vState = 54) and (hState = 571)) or
								((vState = 54) and (hState = 572)) or
								((vState = 54) and (hState = 573)) or
								((vState = 54) and (hState = 574)) or
								((vState = 54) and (hState = 575)) or
								((vState = 54) and (hState = 576)) or
								((vState = 54) and (hState = 579)) or
								((vState = 54) and (hState = 580)) or
								((vState = 54) and (hState = 581)) or
								((vState = 54) and (hState = 582)) or
								((vState = 54) and (hState = 583)) or
								((vState = 54) and (hState = 584)) or
								((vState = 54) and (hState = 585)) or
								((vState = 54) and (hState = 586)) or
								((vState = 54) and (hState = 587)) or
								((vState = 54) and (hState = 595)) or
								((vState = 54) and (hState = 596)) or
								((vState = 54) and (hState = 597)) or
								((vState = 54) and (hState = 598)) or
								((vState = 55) and (hState = 474)) or
								((vState = 55) and (hState = 475)) or
								((vState = 55) and (hState = 481)) or
								((vState = 55) and (hState = 482)) or
								((vState = 55) and (hState = 483)) or
								((vState = 55) and (hState = 484)) or
								((vState = 55) and (hState = 485)) or
								((vState = 55) and (hState = 486)) or
								((vState = 55) and (hState = 487)) or
								((vState = 55) and (hState = 488)) or
								((vState = 55) and (hState = 492)) or
								((vState = 55) and (hState = 493)) or
								((vState = 55) and (hState = 494)) or
								((vState = 55) and (hState = 495)) or
								((vState = 55) and (hState = 496)) or
								((vState = 55) and (hState = 502)) or
								((vState = 55) and (hState = 503)) or
								((vState = 55) and (hState = 504)) or
								((vState = 55) and (hState = 505)) or
								((vState = 55) and (hState = 507)) or
								((vState = 55) and (hState = 508)) or
								((vState = 55) and (hState = 509)) or
								((vState = 55) and (hState = 510)) or
								((vState = 55) and (hState = 512)) or
								((vState = 55) and (hState = 513)) or
								((vState = 55) and (hState = 514)) or
								((vState = 55) and (hState = 515)) or
								((vState = 55) and (hState = 516)) or
								((vState = 55) and (hState = 517)) or
								((vState = 55) and (hState = 518)) or
								((vState = 55) and (hState = 520)) or
								((vState = 55) and (hState = 521)) or
								((vState = 55) and (hState = 522)) or
								((vState = 55) and (hState = 523)) or
								((vState = 55) and (hState = 524)) or
								((vState = 55) and (hState = 525)) or
								((vState = 55) and (hState = 526)) or
								((vState = 55) and (hState = 527)) or
								((vState = 55) and (hState = 528)) or
								((vState = 55) and (hState = 529)) or
								((vState = 55) and (hState = 533)) or
								((vState = 55) and (hState = 534)) or
								((vState = 55) and (hState = 540)) or
								((vState = 55) and (hState = 541)) or
								((vState = 55) and (hState = 542)) or
								((vState = 55) and (hState = 543)) or
								((vState = 55) and (hState = 544)) or
								((vState = 55) and (hState = 554)) or
								((vState = 55) and (hState = 555)) or
								((vState = 55) and (hState = 556)) or
								((vState = 55) and (hState = 561)) or
								((vState = 55) and (hState = 562)) or
								((vState = 55) and (hState = 563)) or
								((vState = 55) and (hState = 564)) or
								((vState = 55) and (hState = 565)) or
								((vState = 55) and (hState = 566)) or
								((vState = 55) and (hState = 567)) or
								((vState = 55) and (hState = 568)) or
								((vState = 55) and (hState = 569)) or
								((vState = 55) and (hState = 570)) or
								((vState = 55) and (hState = 571)) or
								((vState = 55) and (hState = 572)) or
								((vState = 55) and (hState = 573)) or
								((vState = 55) and (hState = 575)) or
								((vState = 55) and (hState = 576)) or
								((vState = 55) and (hState = 580)) or
								((vState = 55) and (hState = 584)) or
								((vState = 55) and (hState = 585)) or
								((vState = 55) and (hState = 586)) or
								((vState = 55) and (hState = 587)) or
								((vState = 55) and (hState = 588)) or
								((vState = 55) and (hState = 597)) or
								((vState = 55) and (hState = 598)) or
								((vState = 55) and (hState = 599)) or
								((vState = 56) and (hState = 474)) or
								((vState = 56) and (hState = 475)) or
								((vState = 56) and (hState = 481)) or
								((vState = 56) and (hState = 482)) or
								((vState = 56) and (hState = 483)) or
								((vState = 56) and (hState = 484)) or
								((vState = 56) and (hState = 485)) or
								((vState = 56) and (hState = 486)) or
								((vState = 56) and (hState = 487)) or
								((vState = 56) and (hState = 488)) or
								((vState = 56) and (hState = 491)) or
								((vState = 56) and (hState = 492)) or
								((vState = 56) and (hState = 493)) or
								((vState = 56) and (hState = 494)) or
								((vState = 56) and (hState = 495)) or
								((vState = 56) and (hState = 496)) or
								((vState = 56) and (hState = 497)) or
								((vState = 56) and (hState = 498)) or
								((vState = 56) and (hState = 501)) or
								((vState = 56) and (hState = 502)) or
								((vState = 56) and (hState = 503)) or
								((vState = 56) and (hState = 504)) or
								((vState = 56) and (hState = 505)) or
								((vState = 56) and (hState = 507)) or
								((vState = 56) and (hState = 508)) or
								((vState = 56) and (hState = 509)) or
								((vState = 56) and (hState = 510)) or
								((vState = 56) and (hState = 512)) or
								((vState = 56) and (hState = 513)) or
								((vState = 56) and (hState = 516)) or
								((vState = 56) and (hState = 517)) or
								((vState = 56) and (hState = 518)) or
								((vState = 56) and (hState = 519)) or
								((vState = 56) and (hState = 520)) or
								((vState = 56) and (hState = 521)) or
								((vState = 56) and (hState = 522)) or
								((vState = 56) and (hState = 523)) or
								((vState = 56) and (hState = 524)) or
								((vState = 56) and (hState = 525)) or
								((vState = 56) and (hState = 526)) or
								((vState = 56) and (hState = 527)) or
								((vState = 56) and (hState = 528)) or
								((vState = 56) and (hState = 529)) or
								((vState = 56) and (hState = 530)) or
								((vState = 56) and (hState = 531)) or
								((vState = 56) and (hState = 533)) or
								((vState = 56) and (hState = 534)) or
								((vState = 56) and (hState = 540)) or
								((vState = 56) and (hState = 541)) or
								((vState = 56) and (hState = 542)) or
								((vState = 56) and (hState = 543)) or
								((vState = 56) and (hState = 544)) or
								((vState = 56) and (hState = 545)) or
								((vState = 56) and (hState = 552)) or
								((vState = 56) and (hState = 553)) or
								((vState = 56) and (hState = 554)) or
								((vState = 56) and (hState = 555)) or
								((vState = 56) and (hState = 560)) or
								((vState = 56) and (hState = 561)) or
								((vState = 56) and (hState = 562)) or
								((vState = 56) and (hState = 563)) or
								((vState = 56) and (hState = 564)) or
								((vState = 56) and (hState = 565)) or
								((vState = 56) and (hState = 566)) or
								((vState = 56) and (hState = 567)) or
								((vState = 56) and (hState = 568)) or
								((vState = 56) and (hState = 569)) or
								((vState = 56) and (hState = 570)) or
								((vState = 56) and (hState = 571)) or
								((vState = 56) and (hState = 572)) or
								((vState = 56) and (hState = 573)) or
								((vState = 56) and (hState = 575)) or
								((vState = 56) and (hState = 576)) or
								((vState = 56) and (hState = 580)) or
								((vState = 56) and (hState = 581)) or
								((vState = 56) and (hState = 586)) or
								((vState = 56) and (hState = 587)) or
								((vState = 56) and (hState = 588)) or
								((vState = 56) and (hState = 589)) or
								((vState = 56) and (hState = 590)) or
								((vState = 56) and (hState = 591)) or
								((vState = 56) and (hState = 597)) or
								((vState = 56) and (hState = 598)) or
								((vState = 56) and (hState = 599)) or
								((vState = 57) and (hState = 473)) or
								((vState = 57) and (hState = 474)) or
								((vState = 57) and (hState = 482)) or
								((vState = 57) and (hState = 483)) or
								((vState = 57) and (hState = 484)) or
								((vState = 57) and (hState = 485)) or
								((vState = 57) and (hState = 486)) or
								((vState = 57) and (hState = 487)) or
								((vState = 57) and (hState = 491)) or
								((vState = 57) and (hState = 492)) or
								((vState = 57) and (hState = 493)) or
								((vState = 57) and (hState = 498)) or
								((vState = 57) and (hState = 499)) or
								((vState = 57) and (hState = 500)) or
								((vState = 57) and (hState = 501)) or
								((vState = 57) and (hState = 502)) or
								((vState = 57) and (hState = 503)) or
								((vState = 57) and (hState = 504)) or
								((vState = 57) and (hState = 507)) or
								((vState = 57) and (hState = 508)) or
								((vState = 57) and (hState = 509)) or
								((vState = 57) and (hState = 510)) or
								((vState = 57) and (hState = 511)) or
								((vState = 57) and (hState = 512)) or
								((vState = 57) and (hState = 517)) or
								((vState = 57) and (hState = 518)) or
								((vState = 57) and (hState = 519)) or
								((vState = 57) and (hState = 520)) or
								((vState = 57) and (hState = 521)) or
								((vState = 57) and (hState = 522)) or
								((vState = 57) and (hState = 523)) or
								((vState = 57) and (hState = 526)) or
								((vState = 57) and (hState = 527)) or
								((vState = 57) and (hState = 528)) or
								((vState = 57) and (hState = 529)) or
								((vState = 57) and (hState = 530)) or
								((vState = 57) and (hState = 531)) or
								((vState = 57) and (hState = 532)) or
								((vState = 57) and (hState = 533)) or
								((vState = 57) and (hState = 534)) or
								((vState = 57) and (hState = 539)) or
								((vState = 57) and (hState = 540)) or
								((vState = 57) and (hState = 541)) or
								((vState = 57) and (hState = 542)) or
								((vState = 57) and (hState = 543)) or
								((vState = 57) and (hState = 544)) or
								((vState = 57) and (hState = 545)) or
								((vState = 57) and (hState = 551)) or
								((vState = 57) and (hState = 552)) or
								((vState = 57) and (hState = 553)) or
								((vState = 57) and (hState = 560)) or
								((vState = 57) and (hState = 561)) or
								((vState = 57) and (hState = 562)) or
								((vState = 57) and (hState = 563)) or
								((vState = 57) and (hState = 564)) or
								((vState = 57) and (hState = 565)) or
								((vState = 57) and (hState = 566)) or
								((vState = 57) and (hState = 567)) or
								((vState = 57) and (hState = 568)) or
								((vState = 57) and (hState = 569)) or
								((vState = 57) and (hState = 570)) or
								((vState = 57) and (hState = 571)) or
								((vState = 57) and (hState = 572)) or
								((vState = 57) and (hState = 573)) or
								((vState = 57) and (hState = 574)) or
								((vState = 57) and (hState = 575)) or
								((vState = 57) and (hState = 576)) or
								((vState = 57) and (hState = 577)) or
								((vState = 57) and (hState = 580)) or
								((vState = 57) and (hState = 581)) or
								((vState = 57) and (hState = 590)) or
								((vState = 57) and (hState = 591)) or
								((vState = 57) and (hState = 592)) or
								((vState = 57) and (hState = 593)) or
								((vState = 57) and (hState = 594)) or
								((vState = 57) and (hState = 595)) or
								((vState = 57) and (hState = 596)) or
								((vState = 57) and (hState = 597)) or
								((vState = 57) and (hState = 598)) or
								((vState = 57) and (hState = 599)) or
								((vState = 58) and (hState = 473)) or
								((vState = 58) and (hState = 474)) or
								((vState = 58) and (hState = 481)) or
								((vState = 58) and (hState = 482)) or
								((vState = 58) and (hState = 483)) or
								((vState = 58) and (hState = 484)) or
								((vState = 58) and (hState = 485)) or
								((vState = 58) and (hState = 486)) or
								((vState = 58) and (hState = 487)) or
								((vState = 58) and (hState = 490)) or
								((vState = 58) and (hState = 491)) or
								((vState = 58) and (hState = 492)) or
								((vState = 58) and (hState = 499)) or
								((vState = 58) and (hState = 500)) or
								((vState = 58) and (hState = 501)) or
								((vState = 58) and (hState = 502)) or
								((vState = 58) and (hState = 503)) or
								((vState = 58) and (hState = 506)) or
								((vState = 58) and (hState = 507)) or
								((vState = 58) and (hState = 508)) or
								((vState = 58) and (hState = 509)) or
								((vState = 58) and (hState = 510)) or
								((vState = 58) and (hState = 511)) or
								((vState = 58) and (hState = 512)) or
								((vState = 58) and (hState = 518)) or
								((vState = 58) and (hState = 519)) or
								((vState = 58) and (hState = 520)) or
								((vState = 58) and (hState = 521)) or
								((vState = 58) and (hState = 527)) or
								((vState = 58) and (hState = 528)) or
								((vState = 58) and (hState = 529)) or
								((vState = 58) and (hState = 530)) or
								((vState = 58) and (hState = 531)) or
								((vState = 58) and (hState = 532)) or
								((vState = 58) and (hState = 533)) or
								((vState = 58) and (hState = 534)) or
								((vState = 58) and (hState = 535)) or
								((vState = 58) and (hState = 538)) or
								((vState = 58) and (hState = 539)) or
								((vState = 58) and (hState = 540)) or
								((vState = 58) and (hState = 543)) or
								((vState = 58) and (hState = 544)) or
								((vState = 58) and (hState = 545)) or
								((vState = 58) and (hState = 546)) or
								((vState = 58) and (hState = 549)) or
								((vState = 58) and (hState = 550)) or
								((vState = 58) and (hState = 551)) or
								((vState = 58) and (hState = 552)) or
								((vState = 58) and (hState = 559)) or
								((vState = 58) and (hState = 560)) or
								((vState = 58) and (hState = 561)) or
								((vState = 58) and (hState = 562)) or
								((vState = 58) and (hState = 563)) or
								((vState = 58) and (hState = 564)) or
								((vState = 58) and (hState = 565)) or
								((vState = 58) and (hState = 566)) or
								((vState = 58) and (hState = 567)) or
								((vState = 58) and (hState = 569)) or
								((vState = 58) and (hState = 570)) or
								((vState = 58) and (hState = 571)) or
								((vState = 58) and (hState = 574)) or
								((vState = 58) and (hState = 575)) or
								((vState = 58) and (hState = 576)) or
								((vState = 58) and (hState = 577)) or
								((vState = 58) and (hState = 580)) or
								((vState = 58) and (hState = 581)) or
								((vState = 58) and (hState = 592)) or
								((vState = 58) and (hState = 593)) or
								((vState = 58) and (hState = 594)) or
								((vState = 58) and (hState = 595)) or
								((vState = 58) and (hState = 596)) or
								((vState = 58) and (hState = 597)) or
								((vState = 59) and (hState = 473)) or
								((vState = 59) and (hState = 474)) or
								((vState = 59) and (hState = 481)) or
								((vState = 59) and (hState = 482)) or
								((vState = 59) and (hState = 483)) or
								((vState = 59) and (hState = 484)) or
								((vState = 59) and (hState = 485)) or
								((vState = 59) and (hState = 486)) or
								((vState = 59) and (hState = 487)) or
								((vState = 59) and (hState = 488)) or
								((vState = 59) and (hState = 489)) or
								((vState = 59) and (hState = 490)) or
								((vState = 59) and (hState = 491)) or
								((vState = 59) and (hState = 500)) or
								((vState = 59) and (hState = 501)) or
								((vState = 59) and (hState = 502)) or
								((vState = 59) and (hState = 503)) or
								((vState = 59) and (hState = 505)) or
								((vState = 59) and (hState = 506)) or
								((vState = 59) and (hState = 507)) or
								((vState = 59) and (hState = 508)) or
								((vState = 59) and (hState = 510)) or
								((vState = 59) and (hState = 511)) or
								((vState = 59) and (hState = 517)) or
								((vState = 59) and (hState = 518)) or
								((vState = 59) and (hState = 519)) or
								((vState = 59) and (hState = 520)) or
								((vState = 59) and (hState = 521)) or
								((vState = 59) and (hState = 527)) or
								((vState = 59) and (hState = 528)) or
								((vState = 59) and (hState = 529)) or
								((vState = 59) and (hState = 531)) or
								((vState = 59) and (hState = 532)) or
								((vState = 59) and (hState = 533)) or
								((vState = 59) and (hState = 534)) or
								((vState = 59) and (hState = 535)) or
								((vState = 59) and (hState = 536)) or
								((vState = 59) and (hState = 537)) or
								((vState = 59) and (hState = 538)) or
								((vState = 59) and (hState = 539)) or
								((vState = 59) and (hState = 540)) or
								((vState = 59) and (hState = 541)) or
								((vState = 59) and (hState = 544)) or
								((vState = 59) and (hState = 545)) or
								((vState = 59) and (hState = 546)) or
								((vState = 59) and (hState = 547)) or
								((vState = 59) and (hState = 548)) or
								((vState = 59) and (hState = 549)) or
								((vState = 59) and (hState = 550)) or
								((vState = 59) and (hState = 558)) or
								((vState = 59) and (hState = 559)) or
								((vState = 59) and (hState = 560)) or
								((vState = 59) and (hState = 561)) or
								((vState = 59) and (hState = 562)) or
								((vState = 59) and (hState = 563)) or
								((vState = 59) and (hState = 564)) or
								((vState = 59) and (hState = 565)) or
								((vState = 59) and (hState = 566)) or
								((vState = 59) and (hState = 569)) or
								((vState = 59) and (hState = 570)) or
								((vState = 59) and (hState = 571)) or
								((vState = 59) and (hState = 572)) or
								((vState = 59) and (hState = 573)) or
								((vState = 59) and (hState = 580)) or
								((vState = 59) and (hState = 581)) or
								((vState = 59) and (hState = 585)) or
								((vState = 59) and (hState = 586)) or
								((vState = 60) and (hState = 473)) or
								((vState = 60) and (hState = 480)) or
								((vState = 60) and (hState = 481)) or
								((vState = 60) and (hState = 482)) or
								((vState = 60) and (hState = 483)) or
								((vState = 60) and (hState = 484)) or
								((vState = 60) and (hState = 485)) or
								((vState = 60) and (hState = 486)) or
								((vState = 60) and (hState = 487)) or
								((vState = 60) and (hState = 488)) or
								((vState = 60) and (hState = 489)) or
								((vState = 60) and (hState = 490)) or
								((vState = 60) and (hState = 491)) or
								((vState = 60) and (hState = 499)) or
								((vState = 60) and (hState = 500)) or
								((vState = 60) and (hState = 501)) or
								((vState = 60) and (hState = 502)) or
								((vState = 60) and (hState = 503)) or
								((vState = 60) and (hState = 504)) or
								((vState = 60) and (hState = 505)) or
								((vState = 60) and (hState = 506)) or
								((vState = 60) and (hState = 507)) or
								((vState = 60) and (hState = 508)) or
								((vState = 60) and (hState = 509)) or
								((vState = 60) and (hState = 510)) or
								((vState = 60) and (hState = 515)) or
								((vState = 60) and (hState = 516)) or
								((vState = 60) and (hState = 517)) or
								((vState = 60) and (hState = 518)) or
								((vState = 60) and (hState = 519)) or
								((vState = 60) and (hState = 520)) or
								((vState = 60) and (hState = 521)) or
								((vState = 60) and (hState = 522)) or
								((vState = 60) and (hState = 527)) or
								((vState = 60) and (hState = 528)) or
								((vState = 60) and (hState = 529)) or
								((vState = 60) and (hState = 533)) or
								((vState = 60) and (hState = 534)) or
								((vState = 60) and (hState = 535)) or
								((vState = 60) and (hState = 536)) or
								((vState = 60) and (hState = 537)) or
								((vState = 60) and (hState = 538)) or
								((vState = 60) and (hState = 539)) or
								((vState = 60) and (hState = 540)) or
								((vState = 60) and (hState = 541)) or
								((vState = 60) and (hState = 545)) or
								((vState = 60) and (hState = 546)) or
								((vState = 60) and (hState = 547)) or
								((vState = 60) and (hState = 548)) or
								((vState = 60) and (hState = 549)) or
								((vState = 60) and (hState = 557)) or
								((vState = 60) and (hState = 558)) or
								((vState = 60) and (hState = 560)) or
								((vState = 60) and (hState = 561)) or
								((vState = 60) and (hState = 562)) or
								((vState = 60) and (hState = 563)) or
								((vState = 60) and (hState = 564)) or
								((vState = 60) and (hState = 565)) or
								((vState = 60) and (hState = 568)) or
								((vState = 60) and (hState = 569)) or
								((vState = 60) and (hState = 571)) or
								((vState = 60) and (hState = 572)) or
								((vState = 60) and (hState = 573)) or
								((vState = 60) and (hState = 574)) or
								((vState = 60) and (hState = 575)) or
								((vState = 60) and (hState = 580)) or
								((vState = 60) and (hState = 581)) or
								((vState = 60) and (hState = 582)) or
								((vState = 60) and (hState = 583)) or
								((vState = 60) and (hState = 584)) or
								((vState = 60) and (hState = 585)) or
								((vState = 60) and (hState = 586)) or
								((vState = 61) and (hState = 472)) or
								((vState = 61) and (hState = 473)) or
								((vState = 61) and (hState = 479)) or
								((vState = 61) and (hState = 480)) or
								((vState = 61) and (hState = 481)) or
								((vState = 61) and (hState = 482)) or
								((vState = 61) and (hState = 483)) or
								((vState = 61) and (hState = 484)) or
								((vState = 61) and (hState = 485)) or
								((vState = 61) and (hState = 486)) or
								((vState = 61) and (hState = 487)) or
								((vState = 61) and (hState = 488)) or
								((vState = 61) and (hState = 489)) or
								((vState = 61) and (hState = 490)) or
								((vState = 61) and (hState = 491)) or
								((vState = 61) and (hState = 492)) or
								((vState = 61) and (hState = 499)) or
								((vState = 61) and (hState = 500)) or
								((vState = 61) and (hState = 501)) or
								((vState = 61) and (hState = 502)) or
								((vState = 61) and (hState = 503)) or
								((vState = 61) and (hState = 504)) or
								((vState = 61) and (hState = 505)) or
								((vState = 61) and (hState = 506)) or
								((vState = 61) and (hState = 507)) or
								((vState = 61) and (hState = 508)) or
								((vState = 61) and (hState = 509)) or
								((vState = 61) and (hState = 510)) or
								((vState = 61) and (hState = 514)) or
								((vState = 61) and (hState = 515)) or
								((vState = 61) and (hState = 516)) or
								((vState = 61) and (hState = 518)) or
								((vState = 61) and (hState = 519)) or
								((vState = 61) and (hState = 520)) or
								((vState = 61) and (hState = 521)) or
								((vState = 61) and (hState = 522)) or
								((vState = 61) and (hState = 523)) or
								((vState = 61) and (hState = 526)) or
								((vState = 61) and (hState = 527)) or
								((vState = 61) and (hState = 528)) or
								((vState = 61) and (hState = 529)) or
								((vState = 61) and (hState = 530)) or
								((vState = 61) and (hState = 533)) or
								((vState = 61) and (hState = 534)) or
								((vState = 61) and (hState = 535)) or
								((vState = 61) and (hState = 536)) or
								((vState = 61) and (hState = 537)) or
								((vState = 61) and (hState = 538)) or
								((vState = 61) and (hState = 539)) or
								((vState = 61) and (hState = 540)) or
								((vState = 61) and (hState = 541)) or
								((vState = 61) and (hState = 546)) or
								((vState = 61) and (hState = 547)) or
								((vState = 61) and (hState = 548)) or
								((vState = 61) and (hState = 549)) or
								((vState = 61) and (hState = 556)) or
								((vState = 61) and (hState = 557)) or
								((vState = 61) and (hState = 561)) or
								((vState = 61) and (hState = 562)) or
								((vState = 61) and (hState = 563)) or
								((vState = 61) and (hState = 564)) or
								((vState = 61) and (hState = 565)) or
								((vState = 61) and (hState = 567)) or
								((vState = 61) and (hState = 568)) or
								((vState = 61) and (hState = 573)) or
								((vState = 61) and (hState = 574)) or
								((vState = 61) and (hState = 575)) or
								((vState = 61) and (hState = 576)) or
								((vState = 61) and (hState = 577)) or
								((vState = 61) and (hState = 579)) or
								((vState = 61) and (hState = 580)) or
								((vState = 61) and (hState = 581)) or
								((vState = 61) and (hState = 582)) or
								((vState = 61) and (hState = 583)) or
								((vState = 61) and (hState = 584)) or
								((vState = 61) and (hState = 585)) or
								((vState = 61) and (hState = 586)) or
								((vState = 62) and (hState = 472)) or
								((vState = 62) and (hState = 473)) or
								((vState = 62) and (hState = 478)) or
								((vState = 62) and (hState = 479)) or
								((vState = 62) and (hState = 480)) or
								((vState = 62) and (hState = 482)) or
								((vState = 62) and (hState = 483)) or
								((vState = 62) and (hState = 484)) or
								((vState = 62) and (hState = 485)) or
								((vState = 62) and (hState = 486)) or
								((vState = 62) and (hState = 487)) or
								((vState = 62) and (hState = 488)) or
								((vState = 62) and (hState = 489)) or
								((vState = 62) and (hState = 490)) or
								((vState = 62) and (hState = 491)) or
								((vState = 62) and (hState = 492)) or
								((vState = 62) and (hState = 493)) or
								((vState = 62) and (hState = 494)) or
								((vState = 62) and (hState = 498)) or
								((vState = 62) and (hState = 499)) or
								((vState = 62) and (hState = 500)) or
								((vState = 62) and (hState = 501)) or
								((vState = 62) and (hState = 502)) or
								((vState = 62) and (hState = 503)) or
								((vState = 62) and (hState = 504)) or
								((vState = 62) and (hState = 505)) or
								((vState = 62) and (hState = 506)) or
								((vState = 62) and (hState = 507)) or
								((vState = 62) and (hState = 508)) or
								((vState = 62) and (hState = 509)) or
								((vState = 62) and (hState = 514)) or
								((vState = 62) and (hState = 515)) or
								((vState = 62) and (hState = 518)) or
								((vState = 62) and (hState = 519)) or
								((vState = 62) and (hState = 521)) or
								((vState = 62) and (hState = 522)) or
								((vState = 62) and (hState = 523)) or
								((vState = 62) and (hState = 524)) or
								((vState = 62) and (hState = 526)) or
								((vState = 62) and (hState = 527)) or
								((vState = 62) and (hState = 529)) or
								((vState = 62) and (hState = 530)) or
								((vState = 62) and (hState = 531)) or
								((vState = 62) and (hState = 533)) or
								((vState = 62) and (hState = 534)) or
								((vState = 62) and (hState = 535)) or
								((vState = 62) and (hState = 536)) or
								((vState = 62) and (hState = 538)) or
								((vState = 62) and (hState = 539)) or
								((vState = 62) and (hState = 540)) or
								((vState = 62) and (hState = 541)) or
								((vState = 62) and (hState = 542)) or
								((vState = 62) and (hState = 543)) or
								((vState = 62) and (hState = 548)) or
								((vState = 62) and (hState = 549)) or
								((vState = 62) and (hState = 555)) or
								((vState = 62) and (hState = 556)) or
								((vState = 62) and (hState = 560)) or
								((vState = 62) and (hState = 561)) or
								((vState = 62) and (hState = 562)) or
								((vState = 62) and (hState = 563)) or
								((vState = 62) and (hState = 564)) or
								((vState = 62) and (hState = 566)) or
								((vState = 62) and (hState = 567)) or
								((vState = 62) and (hState = 568)) or
								((vState = 62) and (hState = 574)) or
								((vState = 62) and (hState = 575)) or
								((vState = 62) and (hState = 576)) or
								((vState = 62) and (hState = 577)) or
								((vState = 62) and (hState = 578)) or
								((vState = 62) and (hState = 579)) or
								((vState = 62) and (hState = 580)) or
								((vState = 62) and (hState = 581)) or
								((vState = 62) and (hState = 582)) or
								((vState = 62) and (hState = 585)) or
								((vState = 62) and (hState = 586)) or
								((vState = 63) and (hState = 472)) or
								((vState = 63) and (hState = 473)) or
								((vState = 63) and (hState = 477)) or
								((vState = 63) and (hState = 478)) or
								((vState = 63) and (hState = 479)) or
								((vState = 63) and (hState = 482)) or
								((vState = 63) and (hState = 483)) or
								((vState = 63) and (hState = 484)) or
								((vState = 63) and (hState = 485)) or
								((vState = 63) and (hState = 486)) or
								((vState = 63) and (hState = 487)) or
								((vState = 63) and (hState = 488)) or
								((vState = 63) and (hState = 489)) or
								((vState = 63) and (hState = 490)) or
								((vState = 63) and (hState = 491)) or
								((vState = 63) and (hState = 492)) or
								((vState = 63) and (hState = 493)) or
								((vState = 63) and (hState = 494)) or
								((vState = 63) and (hState = 498)) or
								((vState = 63) and (hState = 499)) or
								((vState = 63) and (hState = 500)) or
								((vState = 63) and (hState = 501)) or
								((vState = 63) and (hState = 502)) or
								((vState = 63) and (hState = 503)) or
								((vState = 63) and (hState = 504)) or
								((vState = 63) and (hState = 507)) or
								((vState = 63) and (hState = 508)) or
								((vState = 63) and (hState = 509)) or
								((vState = 63) and (hState = 514)) or
								((vState = 63) and (hState = 515)) or
								((vState = 63) and (hState = 518)) or
								((vState = 63) and (hState = 519)) or
								((vState = 63) and (hState = 522)) or
								((vState = 63) and (hState = 523)) or
								((vState = 63) and (hState = 524)) or
								((vState = 63) and (hState = 525)) or
								((vState = 63) and (hState = 526)) or
								((vState = 63) and (hState = 527)) or
								((vState = 63) and (hState = 530)) or
								((vState = 63) and (hState = 531)) or
								((vState = 63) and (hState = 532)) or
								((vState = 63) and (hState = 533)) or
								((vState = 63) and (hState = 534)) or
								((vState = 63) and (hState = 535)) or
								((vState = 63) and (hState = 538)) or
								((vState = 63) and (hState = 539)) or
								((vState = 63) and (hState = 541)) or
								((vState = 63) and (hState = 542)) or
								((vState = 63) and (hState = 543)) or
								((vState = 63) and (hState = 544)) or
								((vState = 63) and (hState = 545)) or
								((vState = 63) and (hState = 549)) or
								((vState = 63) and (hState = 550)) or
								((vState = 63) and (hState = 554)) or
								((vState = 63) and (hState = 555)) or
								((vState = 63) and (hState = 556)) or
								((vState = 63) and (hState = 558)) or
								((vState = 63) and (hState = 559)) or
								((vState = 63) and (hState = 560)) or
								((vState = 63) and (hState = 561)) or
								((vState = 63) and (hState = 562)) or
								((vState = 63) and (hState = 563)) or
								((vState = 63) and (hState = 564)) or
								((vState = 63) and (hState = 565)) or
								((vState = 63) and (hState = 566)) or
								((vState = 63) and (hState = 567)) or
								((vState = 63) and (hState = 573)) or
								((vState = 63) and (hState = 574)) or
								((vState = 63) and (hState = 575)) or
								((vState = 63) and (hState = 576)) or
								((vState = 63) and (hState = 577)) or
								((vState = 63) and (hState = 578)) or
								((vState = 63) and (hState = 579)) or
								((vState = 63) and (hState = 580)) or
								((vState = 63) and (hState = 581)) or
								((vState = 63) and (hState = 582)) or
								((vState = 63) and (hState = 583)) or
								((vState = 63) and (hState = 584)) or
								((vState = 63) and (hState = 585)) or
								((vState = 63) and (hState = 586)) or
								((vState = 63) and (hState = 587)) or
								((vState = 63) and (hState = 588)) or
								((vState = 63) and (hState = 589)) or
								((vState = 63) and (hState = 590)) or
								((vState = 63) and (hState = 591)) or
								((vState = 63) and (hState = 592)) or
								((vState = 63) and (hState = 593)) or
								((vState = 63) and (hState = 594)) or
								((vState = 63) and (hState = 595)) or
								((vState = 63) and (hState = 596)) or
								((vState = 64) and (hState = 471)) or
								((vState = 64) and (hState = 472)) or
								((vState = 64) and (hState = 477)) or
								((vState = 64) and (hState = 478)) or
								((vState = 64) and (hState = 482)) or
								((vState = 64) and (hState = 483)) or
								((vState = 64) and (hState = 484)) or
								((vState = 64) and (hState = 485)) or
								((vState = 64) and (hState = 486)) or
								((vState = 64) and (hState = 487)) or
								((vState = 64) and (hState = 488)) or
								((vState = 64) and (hState = 489)) or
								((vState = 64) and (hState = 490)) or
								((vState = 64) and (hState = 491)) or
								((vState = 64) and (hState = 492)) or
								((vState = 64) and (hState = 493)) or
								((vState = 64) and (hState = 494)) or
								((vState = 64) and (hState = 495)) or
								((vState = 64) and (hState = 496)) or
								((vState = 64) and (hState = 497)) or
								((vState = 64) and (hState = 498)) or
								((vState = 64) and (hState = 499)) or
								((vState = 64) and (hState = 500)) or
								((vState = 64) and (hState = 501)) or
								((vState = 64) and (hState = 502)) or
								((vState = 64) and (hState = 507)) or
								((vState = 64) and (hState = 508)) or
								((vState = 64) and (hState = 514)) or
								((vState = 64) and (hState = 515)) or
								((vState = 64) and (hState = 517)) or
								((vState = 64) and (hState = 518)) or
								((vState = 64) and (hState = 522)) or
								((vState = 64) and (hState = 523)) or
								((vState = 64) and (hState = 524)) or
								((vState = 64) and (hState = 525)) or
								((vState = 64) and (hState = 526)) or
								((vState = 64) and (hState = 527)) or
								((vState = 64) and (hState = 531)) or
								((vState = 64) and (hState = 532)) or
								((vState = 64) and (hState = 533)) or
								((vState = 64) and (hState = 534)) or
								((vState = 64) and (hState = 535)) or
								((vState = 64) and (hState = 538)) or
								((vState = 64) and (hState = 539)) or
								((vState = 64) and (hState = 541)) or
								((vState = 64) and (hState = 544)) or
								((vState = 64) and (hState = 545)) or
								((vState = 64) and (hState = 546)) or
								((vState = 64) and (hState = 547)) or
								((vState = 64) and (hState = 549)) or
								((vState = 64) and (hState = 550)) or
								((vState = 64) and (hState = 551)) or
								((vState = 64) and (hState = 552)) or
								((vState = 64) and (hState = 553)) or
								((vState = 64) and (hState = 554)) or
								((vState = 64) and (hState = 555)) or
								((vState = 64) and (hState = 556)) or
								((vState = 64) and (hState = 557)) or
								((vState = 64) and (hState = 558)) or
								((vState = 64) and (hState = 559)) or
								((vState = 64) and (hState = 560)) or
								((vState = 64) and (hState = 561)) or
								((vState = 64) and (hState = 562)) or
								((vState = 64) and (hState = 563)) or
								((vState = 64) and (hState = 564)) or
								((vState = 64) and (hState = 565)) or
								((vState = 64) and (hState = 566)) or
								((vState = 64) and (hState = 567)) or
								((vState = 64) and (hState = 571)) or
								((vState = 64) and (hState = 572)) or
								((vState = 64) and (hState = 573)) or
								((vState = 64) and (hState = 574)) or
								((vState = 64) and (hState = 575)) or
								((vState = 64) and (hState = 576)) or
								((vState = 64) and (hState = 577)) or
								((vState = 64) and (hState = 578)) or
								((vState = 64) and (hState = 579)) or
								((vState = 64) and (hState = 580)) or
								((vState = 64) and (hState = 581)) or
								((vState = 64) and (hState = 582)) or
								((vState = 64) and (hState = 583)) or
								((vState = 64) and (hState = 584)) or
								((vState = 64) and (hState = 585)) or
								((vState = 64) and (hState = 586)) or
								((vState = 64) and (hState = 587)) or
								((vState = 64) and (hState = 590)) or
								((vState = 64) and (hState = 591)) or
								((vState = 64) and (hState = 592)) or
								((vState = 64) and (hState = 593)) or
								((vState = 64) and (hState = 594)) or
								((vState = 64) and (hState = 595)) or
								((vState = 64) and (hState = 596)) or
								((vState = 65) and (hState = 471)) or
								((vState = 65) and (hState = 472)) or
								((vState = 65) and (hState = 477)) or
								((vState = 65) and (hState = 482)) or
								((vState = 65) and (hState = 483)) or
								((vState = 65) and (hState = 484)) or
								((vState = 65) and (hState = 485)) or
								((vState = 65) and (hState = 486)) or
								((vState = 65) and (hState = 487)) or
								((vState = 65) and (hState = 488)) or
								((vState = 65) and (hState = 494)) or
								((vState = 65) and (hState = 495)) or
								((vState = 65) and (hState = 496)) or
								((vState = 65) and (hState = 497)) or
								((vState = 65) and (hState = 498)) or
								((vState = 65) and (hState = 499)) or
								((vState = 65) and (hState = 500)) or
								((vState = 65) and (hState = 501)) or
								((vState = 65) and (hState = 502)) or
								((vState = 65) and (hState = 503)) or
								((vState = 65) and (hState = 504)) or
								((vState = 65) and (hState = 505)) or
								((vState = 65) and (hState = 506)) or
								((vState = 65) and (hState = 507)) or
								((vState = 65) and (hState = 508)) or
								((vState = 65) and (hState = 509)) or
								((vState = 65) and (hState = 515)) or
								((vState = 65) and (hState = 516)) or
								((vState = 65) and (hState = 517)) or
								((vState = 65) and (hState = 518)) or
								((vState = 65) and (hState = 522)) or
								((vState = 65) and (hState = 523)) or
								((vState = 65) and (hState = 525)) or
								((vState = 65) and (hState = 526)) or
								((vState = 65) and (hState = 527)) or
								((vState = 65) and (hState = 531)) or
								((vState = 65) and (hState = 532)) or
								((vState = 65) and (hState = 533)) or
								((vState = 65) and (hState = 534)) or
								((vState = 65) and (hState = 535)) or
								((vState = 65) and (hState = 536)) or
								((vState = 65) and (hState = 537)) or
								((vState = 65) and (hState = 538)) or
								((vState = 65) and (hState = 539)) or
								((vState = 65) and (hState = 540)) or
								((vState = 65) and (hState = 541)) or
								((vState = 65) and (hState = 544)) or
								((vState = 65) and (hState = 545)) or
								((vState = 65) and (hState = 546)) or
								((vState = 65) and (hState = 547)) or
								((vState = 65) and (hState = 548)) or
								((vState = 65) and (hState = 549)) or
								((vState = 65) and (hState = 550)) or
								((vState = 65) and (hState = 551)) or
								((vState = 65) and (hState = 552)) or
								((vState = 65) and (hState = 553)) or
								((vState = 65) and (hState = 554)) or
								((vState = 65) and (hState = 555)) or
								((vState = 65) and (hState = 556)) or
								((vState = 65) and (hState = 557)) or
								((vState = 65) and (hState = 558)) or
								((vState = 65) and (hState = 559)) or
								((vState = 65) and (hState = 560)) or
								((vState = 65) and (hState = 561)) or
								((vState = 65) and (hState = 562)) or
								((vState = 65) and (hState = 564)) or
								((vState = 65) and (hState = 565)) or
								((vState = 65) and (hState = 566)) or
								((vState = 65) and (hState = 567)) or
								((vState = 65) and (hState = 568)) or
								((vState = 65) and (hState = 569)) or
								((vState = 65) and (hState = 570)) or
								((vState = 65) and (hState = 571)) or
								((vState = 65) and (hState = 572)) or
								((vState = 65) and (hState = 573)) or
								((vState = 65) and (hState = 574)) or
								((vState = 65) and (hState = 575)) or
								((vState = 65) and (hState = 576)) or
								((vState = 65) and (hState = 577)) or
								((vState = 65) and (hState = 578)) or
								((vState = 65) and (hState = 579)) or
								((vState = 65) and (hState = 580)) or
								((vState = 65) and (hState = 581)) or
								((vState = 65) and (hState = 582)) or
								((vState = 65) and (hState = 583)) or
								((vState = 65) and (hState = 584)) or
								((vState = 65) and (hState = 585)) or
								((vState = 65) and (hState = 586)) or
								((vState = 65) and (hState = 595)) or
								((vState = 65) and (hState = 596)) or
								((vState = 66) and (hState = 471)) or
								((vState = 66) and (hState = 472)) or
								((vState = 66) and (hState = 482)) or
								((vState = 66) and (hState = 483)) or
								((vState = 66) and (hState = 484)) or
								((vState = 66) and (hState = 485)) or
								((vState = 66) and (hState = 486)) or
								((vState = 66) and (hState = 487)) or
								((vState = 66) and (hState = 488)) or
								((vState = 66) and (hState = 489)) or
								((vState = 66) and (hState = 495)) or
								((vState = 66) and (hState = 496)) or
								((vState = 66) and (hState = 497)) or
								((vState = 66) and (hState = 498)) or
								((vState = 66) and (hState = 499)) or
								((vState = 66) and (hState = 500)) or
								((vState = 66) and (hState = 504)) or
								((vState = 66) and (hState = 505)) or
								((vState = 66) and (hState = 506)) or
								((vState = 66) and (hState = 507)) or
								((vState = 66) and (hState = 508)) or
								((vState = 66) and (hState = 509)) or
								((vState = 66) and (hState = 510)) or
								((vState = 66) and (hState = 511)) or
								((vState = 66) and (hState = 512)) or
								((vState = 66) and (hState = 515)) or
								((vState = 66) and (hState = 516)) or
								((vState = 66) and (hState = 517)) or
								((vState = 66) and (hState = 518)) or
								((vState = 66) and (hState = 522)) or
								((vState = 66) and (hState = 523)) or
								((vState = 66) and (hState = 524)) or
								((vState = 66) and (hState = 525)) or
								((vState = 66) and (hState = 526)) or
								((vState = 66) and (hState = 527)) or
								((vState = 66) and (hState = 530)) or
								((vState = 66) and (hState = 531)) or
								((vState = 66) and (hState = 532)) or
								((vState = 66) and (hState = 533)) or
								((vState = 66) and (hState = 534)) or
								((vState = 66) and (hState = 535)) or
								((vState = 66) and (hState = 536)) or
								((vState = 66) and (hState = 537)) or
								((vState = 66) and (hState = 538)) or
								((vState = 66) and (hState = 539)) or
								((vState = 66) and (hState = 540)) or
								((vState = 66) and (hState = 541)) or
								((vState = 66) and (hState = 543)) or
								((vState = 66) and (hState = 544)) or
								((vState = 66) and (hState = 545)) or
								((vState = 66) and (hState = 548)) or
								((vState = 66) and (hState = 549)) or
								((vState = 66) and (hState = 550)) or
								((vState = 66) and (hState = 551)) or
								((vState = 66) and (hState = 552)) or
								((vState = 66) and (hState = 553)) or
								((vState = 66) and (hState = 555)) or
								((vState = 66) and (hState = 556)) or
								((vState = 66) and (hState = 557)) or
								((vState = 66) and (hState = 558)) or
								((vState = 66) and (hState = 559)) or
								((vState = 66) and (hState = 560)) or
								((vState = 66) and (hState = 561)) or
								((vState = 66) and (hState = 562)) or
								((vState = 66) and (hState = 563)) or
								((vState = 66) and (hState = 564)) or
								((vState = 66) and (hState = 565)) or
								((vState = 66) and (hState = 566)) or
								((vState = 66) and (hState = 567)) or
								((vState = 66) and (hState = 568)) or
								((vState = 66) and (hState = 569)) or
								((vState = 66) and (hState = 570)) or
								((vState = 66) and (hState = 571)) or
								((vState = 66) and (hState = 572)) or
								((vState = 66) and (hState = 573)) or
								((vState = 66) and (hState = 574)) or
								((vState = 66) and (hState = 576)) or
								((vState = 66) and (hState = 577)) or
								((vState = 66) and (hState = 580)) or
								((vState = 66) and (hState = 581)) or
								((vState = 66) and (hState = 582)) or
								((vState = 66) and (hState = 583)) or
								((vState = 66) and (hState = 584)) or
								((vState = 66) and (hState = 585)) or
								((vState = 66) and (hState = 586)) or
								((vState = 66) and (hState = 587)) or
								((vState = 66) and (hState = 588)) or
								((vState = 66) and (hState = 589)) or
								((vState = 66) and (hState = 595)) or
								((vState = 67) and (hState = 470)) or
								((vState = 67) and (hState = 471)) or
								((vState = 67) and (hState = 482)) or
								((vState = 67) and (hState = 483)) or
								((vState = 67) and (hState = 484)) or
								((vState = 67) and (hState = 485)) or
								((vState = 67) and (hState = 486)) or
								((vState = 67) and (hState = 487)) or
								((vState = 67) and (hState = 488)) or
								((vState = 67) and (hState = 489)) or
								((vState = 67) and (hState = 490)) or
								((vState = 67) and (hState = 491)) or
								((vState = 67) and (hState = 494)) or
								((vState = 67) and (hState = 495)) or
								((vState = 67) and (hState = 496)) or
								((vState = 67) and (hState = 497)) or
								((vState = 67) and (hState = 498)) or
								((vState = 67) and (hState = 499)) or
								((vState = 67) and (hState = 507)) or
								((vState = 67) and (hState = 508)) or
								((vState = 67) and (hState = 511)) or
								((vState = 67) and (hState = 512)) or
								((vState = 67) and (hState = 513)) or
								((vState = 67) and (hState = 515)) or
								((vState = 67) and (hState = 516)) or
								((vState = 67) and (hState = 517)) or
								((vState = 67) and (hState = 522)) or
								((vState = 67) and (hState = 523)) or
								((vState = 67) and (hState = 524)) or
								((vState = 67) and (hState = 525)) or
								((vState = 67) and (hState = 526)) or
								((vState = 67) and (hState = 527)) or
								((vState = 67) and (hState = 528)) or
								((vState = 67) and (hState = 529)) or
								((vState = 67) and (hState = 530)) or
								((vState = 67) and (hState = 531)) or
								((vState = 67) and (hState = 533)) or
								((vState = 67) and (hState = 534)) or
								((vState = 67) and (hState = 537)) or
								((vState = 67) and (hState = 538)) or
								((vState = 67) and (hState = 539)) or
								((vState = 67) and (hState = 540)) or
								((vState = 67) and (hState = 541)) or
								((vState = 67) and (hState = 542)) or
								((vState = 67) and (hState = 543)) or
								((vState = 67) and (hState = 544)) or
								((vState = 67) and (hState = 545)) or
								((vState = 67) and (hState = 550)) or
								((vState = 67) and (hState = 551)) or
								((vState = 67) and (hState = 552)) or
								((vState = 67) and (hState = 553)) or
								((vState = 67) and (hState = 554)) or
								((vState = 67) and (hState = 555)) or
								((vState = 67) and (hState = 556)) or
								((vState = 67) and (hState = 557)) or
								((vState = 67) and (hState = 559)) or
								((vState = 67) and (hState = 560)) or
								((vState = 67) and (hState = 561)) or
								((vState = 67) and (hState = 562)) or
								((vState = 67) and (hState = 563)) or
								((vState = 67) and (hState = 564)) or
								((vState = 67) and (hState = 565)) or
								((vState = 67) and (hState = 566)) or
								((vState = 67) and (hState = 567)) or
								((vState = 67) and (hState = 568)) or
								((vState = 67) and (hState = 569)) or
								((vState = 67) and (hState = 570)) or
								((vState = 67) and (hState = 571)) or
								((vState = 67) and (hState = 572)) or
								((vState = 67) and (hState = 575)) or
								((vState = 67) and (hState = 576)) or
								((vState = 67) and (hState = 577)) or
								((vState = 67) and (hState = 578)) or
								((vState = 67) and (hState = 581)) or
								((vState = 67) and (hState = 582)) or
								((vState = 67) and (hState = 583)) or
								((vState = 67) and (hState = 584)) or
								((vState = 67) and (hState = 585)) or
								((vState = 67) and (hState = 586)) or
								((vState = 67) and (hState = 587)) or
								((vState = 67) and (hState = 588)) or
								((vState = 67) and (hState = 589)) or
								((vState = 67) and (hState = 590)) or
								((vState = 67) and (hState = 591)) or
								((vState = 67) and (hState = 592)) or
								((vState = 67) and (hState = 595)) or
								((vState = 68) and (hState = 470)) or
								((vState = 68) and (hState = 471)) or
								((vState = 68) and (hState = 482)) or
								((vState = 68) and (hState = 483)) or
								((vState = 68) and (hState = 484)) or
								((vState = 68) and (hState = 485)) or
								((vState = 68) and (hState = 486)) or
								((vState = 68) and (hState = 487)) or
								((vState = 68) and (hState = 488)) or
								((vState = 68) and (hState = 489)) or
								((vState = 68) and (hState = 490)) or
								((vState = 68) and (hState = 491)) or
								((vState = 68) and (hState = 492)) or
								((vState = 68) and (hState = 493)) or
								((vState = 68) and (hState = 494)) or
								((vState = 68) and (hState = 495)) or
								((vState = 68) and (hState = 496)) or
								((vState = 68) and (hState = 497)) or
								((vState = 68) and (hState = 498)) or
								((vState = 68) and (hState = 499)) or
								((vState = 68) and (hState = 500)) or
								((vState = 68) and (hState = 507)) or
								((vState = 68) and (hState = 512)) or
								((vState = 68) and (hState = 513)) or
								((vState = 68) and (hState = 516)) or
								((vState = 68) and (hState = 517)) or
								((vState = 68) and (hState = 522)) or
								((vState = 68) and (hState = 523)) or
								((vState = 68) and (hState = 524)) or
								((vState = 68) and (hState = 527)) or
								((vState = 68) and (hState = 528)) or
								((vState = 68) and (hState = 529)) or
								((vState = 68) and (hState = 530)) or
								((vState = 68) and (hState = 533)) or
								((vState = 68) and (hState = 534)) or
								((vState = 68) and (hState = 537)) or
								((vState = 68) and (hState = 538)) or
								((vState = 68) and (hState = 541)) or
								((vState = 68) and (hState = 542)) or
								((vState = 68) and (hState = 543)) or
								((vState = 68) and (hState = 544)) or
								((vState = 68) and (hState = 545)) or
								((vState = 68) and (hState = 546)) or
								((vState = 68) and (hState = 552)) or
								((vState = 68) and (hState = 553)) or
								((vState = 68) and (hState = 554)) or
								((vState = 68) and (hState = 555)) or
								((vState = 68) and (hState = 556)) or
								((vState = 68) and (hState = 560)) or
								((vState = 68) and (hState = 561)) or
								((vState = 68) and (hState = 562)) or
								((vState = 68) and (hState = 563)) or
								((vState = 68) and (hState = 564)) or
								((vState = 68) and (hState = 565)) or
								((vState = 68) and (hState = 566)) or
								((vState = 68) and (hState = 567)) or
								((vState = 68) and (hState = 568)) or
								((vState = 68) and (hState = 569)) or
								((vState = 68) and (hState = 570)) or
								((vState = 68) and (hState = 571)) or
								((vState = 68) and (hState = 575)) or
								((vState = 68) and (hState = 576)) or
								((vState = 68) and (hState = 577)) or
								((vState = 68) and (hState = 578)) or
								((vState = 68) and (hState = 579)) or
								((vState = 68) and (hState = 580)) or
								((vState = 68) and (hState = 581)) or
								((vState = 68) and (hState = 582)) or
								((vState = 68) and (hState = 583)) or
								((vState = 68) and (hState = 584)) or
								((vState = 68) and (hState = 585)) or
								((vState = 68) and (hState = 586)) or
								((vState = 68) and (hState = 587)) or
								((vState = 68) and (hState = 588)) or
								((vState = 68) and (hState = 589)) or
								((vState = 68) and (hState = 590)) or
								((vState = 68) and (hState = 591)) or
								((vState = 68) and (hState = 592)) or
								((vState = 68) and (hState = 593)) or
								((vState = 68) and (hState = 594)) or
								((vState = 68) and (hState = 595)) or
								((vState = 68) and (hState = 596)) or
								((vState = 69) and (hState = 470)) or
								((vState = 69) and (hState = 471)) or
								((vState = 69) and (hState = 481)) or
								((vState = 69) and (hState = 482)) or
								((vState = 69) and (hState = 483)) or
								((vState = 69) and (hState = 484)) or
								((vState = 69) and (hState = 486)) or
								((vState = 69) and (hState = 487)) or
								((vState = 69) and (hState = 488)) or
								((vState = 69) and (hState = 491)) or
								((vState = 69) and (hState = 492)) or
								((vState = 69) and (hState = 493)) or
								((vState = 69) and (hState = 494)) or
								((vState = 69) and (hState = 495)) or
								((vState = 69) and (hState = 496)) or
								((vState = 69) and (hState = 497)) or
								((vState = 69) and (hState = 498)) or
								((vState = 69) and (hState = 499)) or
								((vState = 69) and (hState = 500)) or
								((vState = 69) and (hState = 501)) or
								((vState = 69) and (hState = 502)) or
								((vState = 69) and (hState = 503)) or
								((vState = 69) and (hState = 504)) or
								((vState = 69) and (hState = 506)) or
								((vState = 69) and (hState = 507)) or
								((vState = 69) and (hState = 513)) or
								((vState = 69) and (hState = 514)) or
								((vState = 69) and (hState = 515)) or
								((vState = 69) and (hState = 516)) or
								((vState = 69) and (hState = 517)) or
								((vState = 69) and (hState = 522)) or
								((vState = 69) and (hState = 523)) or
								((vState = 69) and (hState = 524)) or
								((vState = 69) and (hState = 533)) or
								((vState = 69) and (hState = 534)) or
								((vState = 69) and (hState = 535)) or
								((vState = 69) and (hState = 536)) or
								((vState = 69) and (hState = 537)) or
								((vState = 69) and (hState = 538)) or
								((vState = 69) and (hState = 539)) or
								((vState = 69) and (hState = 540)) or
								((vState = 69) and (hState = 541)) or
								((vState = 69) and (hState = 542)) or
								((vState = 69) and (hState = 543)) or
								((vState = 69) and (hState = 544)) or
								((vState = 69) and (hState = 545)) or
								((vState = 69) and (hState = 546)) or
								((vState = 69) and (hState = 547)) or
								((vState = 69) and (hState = 548)) or
								((vState = 69) and (hState = 549)) or
								((vState = 69) and (hState = 553)) or
								((vState = 69) and (hState = 554)) or
								((vState = 69) and (hState = 555)) or
								((vState = 69) and (hState = 556)) or
								((vState = 69) and (hState = 557)) or
								((vState = 69) and (hState = 558)) or
								((vState = 69) and (hState = 559)) or
								((vState = 69) and (hState = 560)) or
								((vState = 69) and (hState = 561)) or
								((vState = 69) and (hState = 562)) or
								((vState = 69) and (hState = 563)) or
								((vState = 69) and (hState = 564)) or
								((vState = 69) and (hState = 565)) or
								((vState = 69) and (hState = 566)) or
								((vState = 69) and (hState = 567)) or
								((vState = 69) and (hState = 568)) or
								((vState = 69) and (hState = 570)) or
								((vState = 69) and (hState = 571)) or
								((vState = 69) and (hState = 572)) or
								((vState = 69) and (hState = 574)) or
								((vState = 69) and (hState = 575)) or
								((vState = 69) and (hState = 576)) or
								((vState = 69) and (hState = 577)) or
								((vState = 69) and (hState = 578)) or
								((vState = 69) and (hState = 579)) or
								((vState = 69) and (hState = 580)) or
								((vState = 69) and (hState = 581)) or
								((vState = 69) and (hState = 582)) or
								((vState = 69) and (hState = 583)) or
								((vState = 69) and (hState = 584)) or
								((vState = 69) and (hState = 585)) or
								((vState = 69) and (hState = 586)) or
								((vState = 69) and (hState = 587)) or
								((vState = 69) and (hState = 588)) or
								((vState = 69) and (hState = 591)) or
								((vState = 69) and (hState = 592)) or
								((vState = 69) and (hState = 593)) or
								((vState = 69) and (hState = 594)) or
								((vState = 69) and (hState = 595)) or
								((vState = 69) and (hState = 596)) or
								((vState = 69) and (hState = 597)) or
								((vState = 70) and (hState = 469)) or
								((vState = 70) and (hState = 470)) or
								((vState = 70) and (hState = 471)) or
								((vState = 70) and (hState = 472)) or
								((vState = 70) and (hState = 481)) or
								((vState = 70) and (hState = 482)) or
								((vState = 70) and (hState = 483)) or
								((vState = 70) and (hState = 486)) or
								((vState = 70) and (hState = 487)) or
								((vState = 70) and (hState = 488)) or
								((vState = 70) and (hState = 489)) or
								((vState = 70) and (hState = 490)) or
								((vState = 70) and (hState = 491)) or
								((vState = 70) and (hState = 492)) or
								((vState = 70) and (hState = 493)) or
								((vState = 70) and (hState = 494)) or
								((vState = 70) and (hState = 495)) or
								((vState = 70) and (hState = 496)) or
								((vState = 70) and (hState = 497)) or
								((vState = 70) and (hState = 498)) or
								((vState = 70) and (hState = 499)) or
								((vState = 70) and (hState = 502)) or
								((vState = 70) and (hState = 503)) or
								((vState = 70) and (hState = 504)) or
								((vState = 70) and (hState = 505)) or
								((vState = 70) and (hState = 506)) or
								((vState = 70) and (hState = 507)) or
								((vState = 70) and (hState = 508)) or
								((vState = 70) and (hState = 509)) or
								((vState = 70) and (hState = 510)) or
								((vState = 70) and (hState = 514)) or
								((vState = 70) and (hState = 515)) or
								((vState = 70) and (hState = 516)) or
								((vState = 70) and (hState = 517)) or
								((vState = 70) and (hState = 522)) or
								((vState = 70) and (hState = 523)) or
								((vState = 70) and (hState = 530)) or
								((vState = 70) and (hState = 531)) or
								((vState = 70) and (hState = 532)) or
								((vState = 70) and (hState = 533)) or
								((vState = 70) and (hState = 534)) or
								((vState = 70) and (hState = 535)) or
								((vState = 70) and (hState = 536)) or
								((vState = 70) and (hState = 537)) or
								((vState = 70) and (hState = 538)) or
								((vState = 70) and (hState = 539)) or
								((vState = 70) and (hState = 540)) or
								((vState = 70) and (hState = 541)) or
								((vState = 70) and (hState = 542)) or
								((vState = 70) and (hState = 543)) or
								((vState = 70) and (hState = 544)) or
								((vState = 70) and (hState = 545)) or
								((vState = 70) and (hState = 546)) or
								((vState = 70) and (hState = 547)) or
								((vState = 70) and (hState = 548)) or
								((vState = 70) and (hState = 549)) or
								((vState = 70) and (hState = 550)) or
								((vState = 70) and (hState = 551)) or
								((vState = 70) and (hState = 552)) or
								((vState = 70) and (hState = 553)) or
								((vState = 70) and (hState = 554)) or
								((vState = 70) and (hState = 557)) or
								((vState = 70) and (hState = 558)) or
								((vState = 70) and (hState = 559)) or
								((vState = 70) and (hState = 560)) or
								((vState = 70) and (hState = 565)) or
								((vState = 70) and (hState = 566)) or
								((vState = 70) and (hState = 567)) or
								((vState = 70) and (hState = 568)) or
								((vState = 70) and (hState = 571)) or
								((vState = 70) and (hState = 572)) or
								((vState = 70) and (hState = 573)) or
								((vState = 70) and (hState = 574)) or
								((vState = 70) and (hState = 575)) or
								((vState = 70) and (hState = 578)) or
								((vState = 70) and (hState = 579)) or
								((vState = 70) and (hState = 580)) or
								((vState = 70) and (hState = 581)) or
								((vState = 70) and (hState = 582)) or
								((vState = 70) and (hState = 583)) or
								((vState = 70) and (hState = 584)) or
								((vState = 70) and (hState = 585)) or
								((vState = 70) and (hState = 587)) or
								((vState = 70) and (hState = 588)) or
								((vState = 70) and (hState = 589)) or
								((vState = 70) and (hState = 594)) or
								((vState = 70) and (hState = 595)) or
								((vState = 70) and (hState = 596)) or
								((vState = 70) and (hState = 597)) or
								((vState = 70) and (hState = 598)) or
								((vState = 70) and (hState = 599)) or
								((vState = 71) and (hState = 469)) or
								((vState = 71) and (hState = 470)) or
								((vState = 71) and (hState = 471)) or
								((vState = 71) and (hState = 472)) or
								((vState = 71) and (hState = 473)) or
								((vState = 71) and (hState = 481)) or
								((vState = 71) and (hState = 482)) or
								((vState = 71) and (hState = 487)) or
								((vState = 71) and (hState = 488)) or
								((vState = 71) and (hState = 489)) or
								((vState = 71) and (hState = 490)) or
								((vState = 71) and (hState = 491)) or
								((vState = 71) and (hState = 492)) or
								((vState = 71) and (hState = 493)) or
								((vState = 71) and (hState = 494)) or
								((vState = 71) and (hState = 495)) or
								((vState = 71) and (hState = 496)) or
								((vState = 71) and (hState = 497)) or
								((vState = 71) and (hState = 498)) or
								((vState = 71) and (hState = 506)) or
								((vState = 71) and (hState = 507)) or
								((vState = 71) and (hState = 508)) or
								((vState = 71) and (hState = 509)) or
								((vState = 71) and (hState = 510)) or
								((vState = 71) and (hState = 511)) or
								((vState = 71) and (hState = 512)) or
								((vState = 71) and (hState = 514)) or
								((vState = 71) and (hState = 515)) or
								((vState = 71) and (hState = 516)) or
								((vState = 71) and (hState = 517)) or
								((vState = 71) and (hState = 518)) or
								((vState = 71) and (hState = 521)) or
								((vState = 71) and (hState = 522)) or
								((vState = 71) and (hState = 527)) or
								((vState = 71) and (hState = 528)) or
								((vState = 71) and (hState = 529)) or
								((vState = 71) and (hState = 530)) or
								((vState = 71) and (hState = 531)) or
								((vState = 71) and (hState = 532)) or
								((vState = 71) and (hState = 533)) or
								((vState = 71) and (hState = 534)) or
								((vState = 71) and (hState = 535)) or
								((vState = 71) and (hState = 536)) or
								((vState = 71) and (hState = 537)) or
								((vState = 71) and (hState = 539)) or
								((vState = 71) and (hState = 540)) or
								((vState = 71) and (hState = 541)) or
								((vState = 71) and (hState = 542)) or
								((vState = 71) and (hState = 545)) or
								((vState = 71) and (hState = 546)) or
								((vState = 71) and (hState = 547)) or
								((vState = 71) and (hState = 548)) or
								((vState = 71) and (hState = 550)) or
								((vState = 71) and (hState = 551)) or
								((vState = 71) and (hState = 552)) or
								((vState = 71) and (hState = 553)) or
								((vState = 71) and (hState = 554)) or
								((vState = 71) and (hState = 558)) or
								((vState = 71) and (hState = 559)) or
								((vState = 71) and (hState = 567)) or
								((vState = 71) and (hState = 568)) or
								((vState = 71) and (hState = 569)) or
								((vState = 71) and (hState = 570)) or
								((vState = 71) and (hState = 572)) or
								((vState = 71) and (hState = 573)) or
								((vState = 71) and (hState = 574)) or
								((vState = 71) and (hState = 580)) or
								((vState = 71) and (hState = 581)) or
								((vState = 71) and (hState = 582)) or
								((vState = 71) and (hState = 583)) or
								((vState = 71) and (hState = 584)) or
								((vState = 71) and (hState = 585)) or
								((vState = 71) and (hState = 588)) or
								((vState = 71) and (hState = 589)) or
								((vState = 71) and (hState = 590)) or
								((vState = 71) and (hState = 594)) or
								((vState = 71) and (hState = 595)) or
								((vState = 71) and (hState = 596)) or
								((vState = 71) and (hState = 597)) or
								((vState = 71) and (hState = 598)) or
								((vState = 71) and (hState = 599)) or
								((vState = 72) and (hState = 468)) or
								((vState = 72) and (hState = 469)) or
								((vState = 72) and (hState = 470)) or
								((vState = 72) and (hState = 471)) or
								((vState = 72) and (hState = 472)) or
								((vState = 72) and (hState = 473)) or
								((vState = 72) and (hState = 480)) or
								((vState = 72) and (hState = 481)) or
								((vState = 72) and (hState = 482)) or
								((vState = 72) and (hState = 486)) or
								((vState = 72) and (hState = 487)) or
								((vState = 72) and (hState = 488)) or
								((vState = 72) and (hState = 489)) or
								((vState = 72) and (hState = 490)) or
								((vState = 72) and (hState = 491)) or
								((vState = 72) and (hState = 494)) or
								((vState = 72) and (hState = 495)) or
								((vState = 72) and (hState = 496)) or
								((vState = 72) and (hState = 497)) or
								((vState = 72) and (hState = 498)) or
								((vState = 72) and (hState = 506)) or
								((vState = 72) and (hState = 507)) or
								((vState = 72) and (hState = 508)) or
								((vState = 72) and (hState = 509)) or
								((vState = 72) and (hState = 510)) or
								((vState = 72) and (hState = 511)) or
								((vState = 72) and (hState = 512)) or
								((vState = 72) and (hState = 515)) or
								((vState = 72) and (hState = 516)) or
								((vState = 72) and (hState = 517)) or
								((vState = 72) and (hState = 518)) or
								((vState = 72) and (hState = 520)) or
								((vState = 72) and (hState = 521)) or
								((vState = 72) and (hState = 522)) or
								((vState = 72) and (hState = 524)) or
								((vState = 72) and (hState = 525)) or
								((vState = 72) and (hState = 526)) or
								((vState = 72) and (hState = 527)) or
								((vState = 72) and (hState = 528)) or
								((vState = 72) and (hState = 529)) or
								((vState = 72) and (hState = 533)) or
								((vState = 72) and (hState = 534)) or
								((vState = 72) and (hState = 535)) or
								((vState = 72) and (hState = 536)) or
								((vState = 72) and (hState = 537)) or
								((vState = 72) and (hState = 538)) or
								((vState = 72) and (hState = 539)) or
								((vState = 72) and (hState = 540)) or
								((vState = 72) and (hState = 541)) or
								((vState = 72) and (hState = 542)) or
								((vState = 72) and (hState = 547)) or
								((vState = 72) and (hState = 548)) or
								((vState = 72) and (hState = 549)) or
								((vState = 72) and (hState = 552)) or
								((vState = 72) and (hState = 553)) or
								((vState = 72) and (hState = 558)) or
								((vState = 72) and (hState = 559)) or
								((vState = 72) and (hState = 569)) or
								((vState = 72) and (hState = 570)) or
								((vState = 72) and (hState = 571)) or
								((vState = 72) and (hState = 572)) or
								((vState = 72) and (hState = 573)) or
								((vState = 72) and (hState = 574)) or
								((vState = 72) and (hState = 575)) or
								((vState = 72) and (hState = 581)) or
								((vState = 72) and (hState = 582)) or
								((vState = 72) and (hState = 583)) or
								((vState = 72) and (hState = 584)) or
								((vState = 72) and (hState = 585)) or
								((vState = 72) and (hState = 586)) or
								((vState = 72) and (hState = 587)) or
								((vState = 72) and (hState = 589)) or
								((vState = 72) and (hState = 590)) or
								((vState = 72) and (hState = 591)) or
								((vState = 72) and (hState = 594)) or
								((vState = 72) and (hState = 595)) or
								((vState = 73) and (hState = 467)) or
								((vState = 73) and (hState = 468)) or
								((vState = 73) and (hState = 469)) or
								((vState = 73) and (hState = 470)) or
								((vState = 73) and (hState = 472)) or
								((vState = 73) and (hState = 473)) or
								((vState = 73) and (hState = 480)) or
								((vState = 73) and (hState = 481)) or
								((vState = 73) and (hState = 485)) or
								((vState = 73) and (hState = 486)) or
								((vState = 73) and (hState = 487)) or
								((vState = 73) and (hState = 488)) or
								((vState = 73) and (hState = 489)) or
								((vState = 73) and (hState = 490)) or
								((vState = 73) and (hState = 494)) or
								((vState = 73) and (hState = 495)) or
								((vState = 73) and (hState = 496)) or
								((vState = 73) and (hState = 497)) or
								((vState = 73) and (hState = 498)) or
								((vState = 73) and (hState = 499)) or
								((vState = 73) and (hState = 500)) or
								((vState = 73) and (hState = 506)) or
								((vState = 73) and (hState = 507)) or
								((vState = 73) and (hState = 508)) or
								((vState = 73) and (hState = 509)) or
								((vState = 73) and (hState = 510)) or
								((vState = 73) and (hState = 515)) or
								((vState = 73) and (hState = 516)) or
								((vState = 73) and (hState = 517)) or
								((vState = 73) and (hState = 518)) or
								((vState = 73) and (hState = 519)) or
								((vState = 73) and (hState = 520)) or
								((vState = 73) and (hState = 521)) or
								((vState = 73) and (hState = 522)) or
								((vState = 73) and (hState = 523)) or
								((vState = 73) and (hState = 524)) or
								((vState = 73) and (hState = 525)) or
								((vState = 73) and (hState = 526)) or
								((vState = 73) and (hState = 533)) or
								((vState = 73) and (hState = 534)) or
								((vState = 73) and (hState = 535)) or
								((vState = 73) and (hState = 536)) or
								((vState = 73) and (hState = 537)) or
								((vState = 73) and (hState = 538)) or
								((vState = 73) and (hState = 539)) or
								((vState = 73) and (hState = 541)) or
								((vState = 73) and (hState = 542)) or
								((vState = 73) and (hState = 548)) or
								((vState = 73) and (hState = 549)) or
								((vState = 73) and (hState = 550)) or
								((vState = 73) and (hState = 551)) or
								((vState = 73) and (hState = 552)) or
								((vState = 73) and (hState = 557)) or
								((vState = 73) and (hState = 558)) or
								((vState = 73) and (hState = 566)) or
								((vState = 73) and (hState = 571)) or
								((vState = 73) and (hState = 572)) or
								((vState = 73) and (hState = 573)) or
								((vState = 73) and (hState = 574)) or
								((vState = 73) and (hState = 575)) or
								((vState = 73) and (hState = 576)) or
								((vState = 73) and (hState = 582)) or
								((vState = 73) and (hState = 583)) or
								((vState = 73) and (hState = 584)) or
								((vState = 73) and (hState = 585)) or
								((vState = 73) and (hState = 586)) or
								((vState = 73) and (hState = 587)) or
								((vState = 73) and (hState = 588)) or
								((vState = 73) and (hState = 589)) or
								((vState = 73) and (hState = 590)) or
								((vState = 73) and (hState = 591)) or
								((vState = 73) and (hState = 592)) or
								((vState = 73) and (hState = 593)) or
								((vState = 73) and (hState = 594)) or
								((vState = 73) and (hState = 595)) or
								((vState = 73) and (hState = 599)) or
								((vState = 74) and (hState = 465)) or
								((vState = 74) and (hState = 466)) or
								((vState = 74) and (hState = 467)) or
								((vState = 74) and (hState = 468)) or
								((vState = 74) and (hState = 469)) or
								((vState = 74) and (hState = 472)) or
								((vState = 74) and (hState = 473)) or
								((vState = 74) and (hState = 480)) or
								((vState = 74) and (hState = 481)) or
								((vState = 74) and (hState = 484)) or
								((vState = 74) and (hState = 485)) or
								((vState = 74) and (hState = 486)) or
								((vState = 74) and (hState = 487)) or
								((vState = 74) and (hState = 488)) or
								((vState = 74) and (hState = 489)) or
								((vState = 74) and (hState = 490)) or
								((vState = 74) and (hState = 491)) or
								((vState = 74) and (hState = 493)) or
								((vState = 74) and (hState = 494)) or
								((vState = 74) and (hState = 495)) or
								((vState = 74) and (hState = 496)) or
								((vState = 74) and (hState = 497)) or
								((vState = 74) and (hState = 498)) or
								((vState = 74) and (hState = 499)) or
								((vState = 74) and (hState = 500)) or
								((vState = 74) and (hState = 501)) or
								((vState = 74) and (hState = 505)) or
								((vState = 74) and (hState = 506)) or
								((vState = 74) and (hState = 507)) or
								((vState = 74) and (hState = 508)) or
								((vState = 74) and (hState = 515)) or
								((vState = 74) and (hState = 517)) or
								((vState = 74) and (hState = 518)) or
								((vState = 74) and (hState = 519)) or
								((vState = 74) and (hState = 520)) or
								((vState = 74) and (hState = 521)) or
								((vState = 74) and (hState = 522)) or
								((vState = 74) and (hState = 523)) or
								((vState = 74) and (hState = 534)) or
								((vState = 74) and (hState = 535)) or
								((vState = 74) and (hState = 536)) or
								((vState = 74) and (hState = 537)) or
								((vState = 74) and (hState = 538)) or
								((vState = 74) and (hState = 541)) or
								((vState = 74) and (hState = 542)) or
								((vState = 74) and (hState = 550)) or
								((vState = 74) and (hState = 551)) or
								((vState = 74) and (hState = 552)) or
								((vState = 74) and (hState = 557)) or
								((vState = 74) and (hState = 558)) or
								((vState = 74) and (hState = 565)) or
								((vState = 74) and (hState = 566)) or
								((vState = 74) and (hState = 567)) or
								((vState = 74) and (hState = 575)) or
								((vState = 74) and (hState = 576)) or
								((vState = 74) and (hState = 577)) or
								((vState = 74) and (hState = 583)) or
								((vState = 74) and (hState = 584)) or
								((vState = 74) and (hState = 585)) or
								((vState = 74) and (hState = 586)) or
								((vState = 74) and (hState = 587)) or
								((vState = 74) and (hState = 588)) or
								((vState = 74) and (hState = 589)) or
								((vState = 74) and (hState = 590)) or
								((vState = 74) and (hState = 591)) or
								((vState = 74) and (hState = 592)) or
								((vState = 74) and (hState = 593)) or
								((vState = 74) and (hState = 594)) or
								((vState = 74) and (hState = 595)) or
								((vState = 74) and (hState = 598)) or
								((vState = 74) and (hState = 599)) or
								((vState = 75) and (hState = 464)) or
								((vState = 75) and (hState = 465)) or
								((vState = 75) and (hState = 466)) or
								((vState = 75) and (hState = 468)) or
								((vState = 75) and (hState = 469)) or
								((vState = 75) and (hState = 470)) or
								((vState = 75) and (hState = 471)) or
								((vState = 75) and (hState = 472)) or
								((vState = 75) and (hState = 473)) or
								((vState = 75) and (hState = 480)) or
								((vState = 75) and (hState = 481)) or
								((vState = 75) and (hState = 482)) or
								((vState = 75) and (hState = 483)) or
								((vState = 75) and (hState = 484)) or
								((vState = 75) and (hState = 485)) or
								((vState = 75) and (hState = 486)) or
								((vState = 75) and (hState = 487)) or
								((vState = 75) and (hState = 488)) or
								((vState = 75) and (hState = 489)) or
								((vState = 75) and (hState = 490)) or
								((vState = 75) and (hState = 491)) or
								((vState = 75) and (hState = 492)) or
								((vState = 75) and (hState = 493)) or
								((vState = 75) and (hState = 494)) or
								((vState = 75) and (hState = 495)) or
								((vState = 75) and (hState = 496)) or
								((vState = 75) and (hState = 497)) or
								((vState = 75) and (hState = 498)) or
								((vState = 75) and (hState = 499)) or
								((vState = 75) and (hState = 500)) or
								((vState = 75) and (hState = 501)) or
								((vState = 75) and (hState = 502)) or
								((vState = 75) and (hState = 503)) or
								((vState = 75) and (hState = 504)) or
								((vState = 75) and (hState = 505)) or
								((vState = 75) and (hState = 506)) or
								((vState = 75) and (hState = 514)) or
								((vState = 75) and (hState = 515)) or
								((vState = 75) and (hState = 517)) or
								((vState = 75) and (hState = 518)) or
								((vState = 75) and (hState = 519)) or
								((vState = 75) and (hState = 520)) or
								((vState = 75) and (hState = 535)) or
								((vState = 75) and (hState = 536)) or
								((vState = 75) and (hState = 537)) or
								((vState = 75) and (hState = 538)) or
								((vState = 75) and (hState = 539)) or
								((vState = 75) and (hState = 540)) or
								((vState = 75) and (hState = 541)) or
								((vState = 75) and (hState = 542)) or
								((vState = 75) and (hState = 550)) or
								((vState = 75) and (hState = 551)) or
								((vState = 75) and (hState = 552)) or
								((vState = 75) and (hState = 553)) or
								((vState = 75) and (hState = 556)) or
								((vState = 75) and (hState = 557)) or
								((vState = 75) and (hState = 558)) or
								((vState = 75) and (hState = 559)) or
								((vState = 75) and (hState = 560)) or
								((vState = 75) and (hState = 561)) or
								((vState = 75) and (hState = 565)) or
								((vState = 75) and (hState = 566)) or
								((vState = 75) and (hState = 567)) or
								((vState = 75) and (hState = 568)) or
								((vState = 75) and (hState = 569)) or
								((vState = 75) and (hState = 577)) or
								((vState = 75) and (hState = 578)) or
								((vState = 75) and (hState = 583)) or
								((vState = 75) and (hState = 584)) or
								((vState = 75) and (hState = 585)) or
								((vState = 75) and (hState = 586)) or
								((vState = 75) and (hState = 587)) or
								((vState = 75) and (hState = 588)) or
								((vState = 75) and (hState = 589)) or
								((vState = 75) and (hState = 590)) or
								((vState = 75) and (hState = 591)) or
								((vState = 75) and (hState = 592)) or
								((vState = 75) and (hState = 593)) or
								((vState = 75) and (hState = 594)) or
								((vState = 75) and (hState = 595)) or
								((vState = 75) and (hState = 598)) or
								((vState = 75) and (hState = 599)) or
								((vState = 76) and (hState = 462)) or
								((vState = 76) and (hState = 463)) or
								((vState = 76) and (hState = 464)) or
								((vState = 76) and (hState = 465)) or
								((vState = 76) and (hState = 467)) or
								((vState = 76) and (hState = 468)) or
								((vState = 76) and (hState = 469)) or
								((vState = 76) and (hState = 470)) or
								((vState = 76) and (hState = 471)) or
								((vState = 76) and (hState = 472)) or
								((vState = 76) and (hState = 473)) or
								((vState = 76) and (hState = 480)) or
								((vState = 76) and (hState = 481)) or
								((vState = 76) and (hState = 482)) or
								((vState = 76) and (hState = 483)) or
								((vState = 76) and (hState = 484)) or
								((vState = 76) and (hState = 485)) or
								((vState = 76) and (hState = 486)) or
								((vState = 76) and (hState = 487)) or
								((vState = 76) and (hState = 488)) or
								((vState = 76) and (hState = 489)) or
								((vState = 76) and (hState = 490)) or
								((vState = 76) and (hState = 491)) or
								((vState = 76) and (hState = 492)) or
								((vState = 76) and (hState = 496)) or
								((vState = 76) and (hState = 497)) or
								((vState = 76) and (hState = 498)) or
								((vState = 76) and (hState = 499)) or
								((vState = 76) and (hState = 500)) or
								((vState = 76) and (hState = 501)) or
								((vState = 76) and (hState = 502)) or
								((vState = 76) and (hState = 503)) or
								((vState = 76) and (hState = 504)) or
								((vState = 76) and (hState = 505)) or
								((vState = 76) and (hState = 506)) or
								((vState = 76) and (hState = 514)) or
								((vState = 76) and (hState = 515)) or
								((vState = 76) and (hState = 517)) or
								((vState = 76) and (hState = 518)) or
								((vState = 76) and (hState = 519)) or
								((vState = 76) and (hState = 520)) or
								((vState = 76) and (hState = 534)) or
								((vState = 76) and (hState = 535)) or
								((vState = 76) and (hState = 536)) or
								((vState = 76) and (hState = 539)) or
								((vState = 76) and (hState = 540)) or
								((vState = 76) and (hState = 541)) or
								((vState = 76) and (hState = 542)) or
								((vState = 76) and (hState = 543)) or
								((vState = 76) and (hState = 550)) or
								((vState = 76) and (hState = 551)) or
								((vState = 76) and (hState = 552)) or
								((vState = 76) and (hState = 553)) or
								((vState = 76) and (hState = 554)) or
								((vState = 76) and (hState = 555)) or
								((vState = 76) and (hState = 556)) or
								((vState = 76) and (hState = 557)) or
								((vState = 76) and (hState = 558)) or
								((vState = 76) and (hState = 560)) or
								((vState = 76) and (hState = 561)) or
								((vState = 76) and (hState = 562)) or
								((vState = 76) and (hState = 566)) or
								((vState = 76) and (hState = 567)) or
								((vState = 76) and (hState = 568)) or
								((vState = 76) and (hState = 569)) or
								((vState = 76) and (hState = 570)) or
								((vState = 76) and (hState = 571)) or
								((vState = 76) and (hState = 577)) or
								((vState = 76) and (hState = 578)) or
								((vState = 76) and (hState = 584)) or
								((vState = 76) and (hState = 585)) or
								((vState = 76) and (hState = 586)) or
								((vState = 76) and (hState = 587)) or
								((vState = 76) and (hState = 588)) or
								((vState = 76) and (hState = 589)) or
								((vState = 76) and (hState = 590)) or
								((vState = 76) and (hState = 591)) or
								((vState = 76) and (hState = 592)) or
								((vState = 76) and (hState = 593)) or
								((vState = 76) and (hState = 594)) or
								((vState = 76) and (hState = 595)) or
								((vState = 76) and (hState = 596)) or
								((vState = 76) and (hState = 597)) or
								((vState = 76) and (hState = 598)) or
								((vState = 77) and (hState = 460)) or
								((vState = 77) and (hState = 461)) or
								((vState = 77) and (hState = 462)) or
								((vState = 77) and (hState = 463)) or
								((vState = 77) and (hState = 464)) or
								((vState = 77) and (hState = 465)) or
								((vState = 77) and (hState = 466)) or
								((vState = 77) and (hState = 467)) or
								((vState = 77) and (hState = 468)) or
								((vState = 77) and (hState = 469)) or
								((vState = 77) and (hState = 471)) or
								((vState = 77) and (hState = 472)) or
								((vState = 77) and (hState = 473)) or
								((vState = 77) and (hState = 479)) or
								((vState = 77) and (hState = 480)) or
								((vState = 77) and (hState = 481)) or
								((vState = 77) and (hState = 482)) or
								((vState = 77) and (hState = 483)) or
								((vState = 77) and (hState = 484)) or
								((vState = 77) and (hState = 485)) or
								((vState = 77) and (hState = 486)) or
								((vState = 77) and (hState = 487)) or
								((vState = 77) and (hState = 491)) or
								((vState = 77) and (hState = 492)) or
								((vState = 77) and (hState = 493)) or
								((vState = 77) and (hState = 496)) or
								((vState = 77) and (hState = 497)) or
								((vState = 77) and (hState = 498)) or
								((vState = 77) and (hState = 499)) or
								((vState = 77) and (hState = 500)) or
								((vState = 77) and (hState = 501)) or
								((vState = 77) and (hState = 502)) or
								((vState = 77) and (hState = 503)) or
								((vState = 77) and (hState = 504)) or
								((vState = 77) and (hState = 505)) or
								((vState = 77) and (hState = 506)) or
								((vState = 77) and (hState = 507)) or
								((vState = 77) and (hState = 508)) or
								((vState = 77) and (hState = 509)) or
								((vState = 77) and (hState = 510)) or
								((vState = 77) and (hState = 511)) or
								((vState = 77) and (hState = 512)) or
								((vState = 77) and (hState = 513)) or
								((vState = 77) and (hState = 514)) or
								((vState = 77) and (hState = 515)) or
								((vState = 77) and (hState = 516)) or
								((vState = 77) and (hState = 517)) or
								((vState = 77) and (hState = 518)) or
								((vState = 77) and (hState = 519)) or
								((vState = 77) and (hState = 520)) or
								((vState = 77) and (hState = 521)) or
								((vState = 77) and (hState = 534)) or
								((vState = 77) and (hState = 535)) or
								((vState = 77) and (hState = 536)) or
								((vState = 77) and (hState = 541)) or
								((vState = 77) and (hState = 542)) or
								((vState = 77) and (hState = 543)) or
								((vState = 77) and (hState = 544)) or
								((vState = 77) and (hState = 545)) or
								((vState = 77) and (hState = 546)) or
								((vState = 77) and (hState = 547)) or
								((vState = 77) and (hState = 550)) or
								((vState = 77) and (hState = 551)) or
								((vState = 77) and (hState = 552)) or
								((vState = 77) and (hState = 553)) or
								((vState = 77) and (hState = 554)) or
								((vState = 77) and (hState = 555)) or
								((vState = 77) and (hState = 556)) or
								((vState = 77) and (hState = 561)) or
								((vState = 77) and (hState = 562)) or
								((vState = 77) and (hState = 563)) or
								((vState = 77) and (hState = 566)) or
								((vState = 77) and (hState = 567)) or
								((vState = 77) and (hState = 570)) or
								((vState = 77) and (hState = 571)) or
								((vState = 77) and (hState = 572)) or
								((vState = 77) and (hState = 577)) or
								((vState = 77) and (hState = 578)) or
								((vState = 77) and (hState = 585)) or
								((vState = 77) and (hState = 586)) or
								((vState = 77) and (hState = 587)) or
								((vState = 77) and (hState = 588)) or
								((vState = 77) and (hState = 589)) or
								((vState = 77) and (hState = 590)) or
								((vState = 77) and (hState = 591)) or
								((vState = 77) and (hState = 593)) or
								((vState = 77) and (hState = 594)) or
								((vState = 77) and (hState = 595)) or
								((vState = 77) and (hState = 596)) or
								((vState = 77) and (hState = 597)) or
								((vState = 78) and (hState = 459)) or
								((vState = 78) and (hState = 460)) or
								((vState = 78) and (hState = 461)) or
								((vState = 78) and (hState = 462)) or
								((vState = 78) and (hState = 463)) or
								((vState = 78) and (hState = 464)) or
								((vState = 78) and (hState = 465)) or
								((vState = 78) and (hState = 466)) or
								((vState = 78) and (hState = 467)) or
								((vState = 78) and (hState = 468)) or
								((vState = 78) and (hState = 472)) or
								((vState = 78) and (hState = 473)) or
								((vState = 78) and (hState = 474)) or
								((vState = 78) and (hState = 478)) or
								((vState = 78) and (hState = 479)) or
								((vState = 78) and (hState = 480)) or
								((vState = 78) and (hState = 485)) or
								((vState = 78) and (hState = 486)) or
								((vState = 78) and (hState = 491)) or
								((vState = 78) and (hState = 492)) or
								((vState = 78) and (hState = 493)) or
								((vState = 78) and (hState = 494)) or
								((vState = 78) and (hState = 495)) or
								((vState = 78) and (hState = 496)) or
								((vState = 78) and (hState = 497)) or
								((vState = 78) and (hState = 498)) or
								((vState = 78) and (hState = 499)) or
								((vState = 78) and (hState = 500)) or
								((vState = 78) and (hState = 501)) or
								((vState = 78) and (hState = 502)) or
								((vState = 78) and (hState = 503)) or
								((vState = 78) and (hState = 504)) or
								((vState = 78) and (hState = 505)) or
								((vState = 78) and (hState = 506)) or
								((vState = 78) and (hState = 507)) or
								((vState = 78) and (hState = 508)) or
								((vState = 78) and (hState = 509)) or
								((vState = 78) and (hState = 510)) or
								((vState = 78) and (hState = 511)) or
								((vState = 78) and (hState = 512)) or
								((vState = 78) and (hState = 513)) or
								((vState = 78) and (hState = 514)) or
								((vState = 78) and (hState = 515)) or
								((vState = 78) and (hState = 516)) or
								((vState = 78) and (hState = 517)) or
								((vState = 78) and (hState = 518)) or
								((vState = 78) and (hState = 519)) or
								((vState = 78) and (hState = 520)) or
								((vState = 78) and (hState = 521)) or
								((vState = 78) and (hState = 522)) or
								((vState = 78) and (hState = 524)) or
								((vState = 78) and (hState = 525)) or
								((vState = 78) and (hState = 533)) or
								((vState = 78) and (hState = 534)) or
								((vState = 78) and (hState = 535)) or
								((vState = 78) and (hState = 542)) or
								((vState = 78) and (hState = 543)) or
								((vState = 78) and (hState = 544)) or
								((vState = 78) and (hState = 545)) or
								((vState = 78) and (hState = 546)) or
								((vState = 78) and (hState = 547)) or
								((vState = 78) and (hState = 548)) or
								((vState = 78) and (hState = 549)) or
								((vState = 78) and (hState = 550)) or
								((vState = 78) and (hState = 551)) or
								((vState = 78) and (hState = 552)) or
								((vState = 78) and (hState = 553)) or
								((vState = 78) and (hState = 554)) or
								((vState = 78) and (hState = 555)) or
								((vState = 78) and (hState = 556)) or
								((vState = 78) and (hState = 562)) or
								((vState = 78) and (hState = 563)) or
								((vState = 78) and (hState = 564)) or
								((vState = 78) and (hState = 566)) or
								((vState = 78) and (hState = 567)) or
								((vState = 78) and (hState = 571)) or
								((vState = 78) and (hState = 572)) or
								((vState = 78) and (hState = 573)) or
								((vState = 78) and (hState = 577)) or
								((vState = 78) and (hState = 586)) or
								((vState = 78) and (hState = 587)) or
								((vState = 78) and (hState = 588)) or
								((vState = 78) and (hState = 589)) or
								((vState = 78) and (hState = 590)) or
								((vState = 78) and (hState = 591)) or
								((vState = 78) and (hState = 592)) or
								((vState = 78) and (hState = 593)) or
								((vState = 78) and (hState = 594)) or
								((vState = 78) and (hState = 595)) or
								((vState = 78) and (hState = 596)) or
								((vState = 78) and (hState = 597)) or
								((vState = 78) and (hState = 598)) or
								((vState = 79) and (hState = 457)) or
								((vState = 79) and (hState = 458)) or
								((vState = 79) and (hState = 459)) or
								((vState = 79) and (hState = 460)) or
								((vState = 79) and (hState = 461)) or
								((vState = 79) and (hState = 462)) or
								((vState = 79) and (hState = 463)) or
								((vState = 79) and (hState = 467)) or
								((vState = 79) and (hState = 468)) or
								((vState = 79) and (hState = 472)) or
								((vState = 79) and (hState = 473)) or
								((vState = 79) and (hState = 474)) or
								((vState = 79) and (hState = 475)) or
								((vState = 79) and (hState = 476)) or
								((vState = 79) and (hState = 477)) or
								((vState = 79) and (hState = 478)) or
								((vState = 79) and (hState = 479)) or
								((vState = 79) and (hState = 485)) or
								((vState = 79) and (hState = 486)) or
								((vState = 79) and (hState = 492)) or
								((vState = 79) and (hState = 493)) or
								((vState = 79) and (hState = 494)) or
								((vState = 79) and (hState = 495)) or
								((vState = 79) and (hState = 496)) or
								((vState = 79) and (hState = 497)) or
								((vState = 79) and (hState = 498)) or
								((vState = 79) and (hState = 499)) or
								((vState = 79) and (hState = 500)) or
								((vState = 79) and (hState = 501)) or
								((vState = 79) and (hState = 505)) or
								((vState = 79) and (hState = 506)) or
								((vState = 79) and (hState = 507)) or
								((vState = 79) and (hState = 508)) or
								((vState = 79) and (hState = 509)) or
								((vState = 79) and (hState = 515)) or
								((vState = 79) and (hState = 516)) or
								((vState = 79) and (hState = 517)) or
								((vState = 79) and (hState = 518)) or
								((vState = 79) and (hState = 519)) or
								((vState = 79) and (hState = 520)) or
								((vState = 79) and (hState = 522)) or
								((vState = 79) and (hState = 523)) or
								((vState = 79) and (hState = 524)) or
								((vState = 79) and (hState = 525)) or
								((vState = 79) and (hState = 526)) or
								((vState = 79) and (hState = 533)) or
								((vState = 79) and (hState = 534)) or
								((vState = 79) and (hState = 543)) or
								((vState = 79) and (hState = 544)) or
								((vState = 79) and (hState = 547)) or
								((vState = 79) and (hState = 548)) or
								((vState = 79) and (hState = 549)) or
								((vState = 79) and (hState = 550)) or
								((vState = 79) and (hState = 551)) or
								((vState = 79) and (hState = 552)) or
								((vState = 79) and (hState = 553)) or
								((vState = 79) and (hState = 554)) or
								((vState = 79) and (hState = 555)) or
								((vState = 79) and (hState = 556)) or
								((vState = 79) and (hState = 557)) or
								((vState = 79) and (hState = 558)) or
								((vState = 79) and (hState = 564)) or
								((vState = 79) and (hState = 565)) or
								((vState = 79) and (hState = 567)) or
								((vState = 79) and (hState = 572)) or
								((vState = 79) and (hState = 573)) or
								((vState = 79) and (hState = 574)) or
								((vState = 79) and (hState = 577)) or
								((vState = 79) and (hState = 587)) or
								((vState = 79) and (hState = 588)) or
								((vState = 79) and (hState = 591)) or
								((vState = 79) and (hState = 592)) or
								((vState = 79) and (hState = 593)) or
								((vState = 79) and (hState = 594)) or
								((vState = 79) and (hState = 595)) or
								((vState = 79) and (hState = 596)) or
								((vState = 79) and (hState = 598)) or
								((vState = 80) and (hState = 455)) or
								((vState = 80) and (hState = 456)) or
								((vState = 80) and (hState = 457)) or
								((vState = 80) and (hState = 458)) or
								((vState = 80) and (hState = 459)) or
								((vState = 80) and (hState = 460)) or
								((vState = 80) and (hState = 466)) or
								((vState = 80) and (hState = 467)) or
								((vState = 80) and (hState = 473)) or
								((vState = 80) and (hState = 474)) or
								((vState = 80) and (hState = 475)) or
								((vState = 80) and (hState = 476)) or
								((vState = 80) and (hState = 477)) or
								((vState = 80) and (hState = 485)) or
								((vState = 80) and (hState = 486)) or
								((vState = 80) and (hState = 491)) or
								((vState = 80) and (hState = 492)) or
								((vState = 80) and (hState = 493)) or
								((vState = 80) and (hState = 494)) or
								((vState = 80) and (hState = 495)) or
								((vState = 80) and (hState = 496)) or
								((vState = 80) and (hState = 497)) or
								((vState = 80) and (hState = 498)) or
								((vState = 80) and (hState = 499)) or
								((vState = 80) and (hState = 500)) or
								((vState = 80) and (hState = 501)) or
								((vState = 80) and (hState = 505)) or
								((vState = 80) and (hState = 506)) or
								((vState = 80) and (hState = 507)) or
								((vState = 80) and (hState = 508)) or
								((vState = 80) and (hState = 509)) or
								((vState = 80) and (hState = 510)) or
								((vState = 80) and (hState = 514)) or
								((vState = 80) and (hState = 515)) or
								((vState = 80) and (hState = 516)) or
								((vState = 80) and (hState = 517)) or
								((vState = 80) and (hState = 518)) or
								((vState = 80) and (hState = 519)) or
								((vState = 80) and (hState = 520)) or
								((vState = 80) and (hState = 522)) or
								((vState = 80) and (hState = 523)) or
								((vState = 80) and (hState = 524)) or
								((vState = 80) and (hState = 525)) or
								((vState = 80) and (hState = 526)) or
								((vState = 80) and (hState = 533)) or
								((vState = 80) and (hState = 534)) or
								((vState = 80) and (hState = 544)) or
								((vState = 80) and (hState = 545)) or
								((vState = 80) and (hState = 546)) or
								((vState = 80) and (hState = 547)) or
								((vState = 80) and (hState = 548)) or
								((vState = 80) and (hState = 549)) or
								((vState = 80) and (hState = 550)) or
								((vState = 80) and (hState = 551)) or
								((vState = 80) and (hState = 552)) or
								((vState = 80) and (hState = 553)) or
								((vState = 80) and (hState = 554)) or
								((vState = 80) and (hState = 555)) or
								((vState = 80) and (hState = 556)) or
								((vState = 80) and (hState = 557)) or
								((vState = 80) and (hState = 558)) or
								((vState = 80) and (hState = 559)) or
								((vState = 80) and (hState = 560)) or
								((vState = 80) and (hState = 564)) or
								((vState = 80) and (hState = 565)) or
								((vState = 80) and (hState = 566)) or
								((vState = 80) and (hState = 567)) or
								((vState = 80) and (hState = 572)) or
								((vState = 80) and (hState = 573)) or
								((vState = 80) and (hState = 577)) or
								((vState = 80) and (hState = 582)) or
								((vState = 80) and (hState = 587)) or
								((vState = 80) and (hState = 588)) or
								((vState = 80) and (hState = 589)) or
								((vState = 80) and (hState = 592)) or
								((vState = 80) and (hState = 593)) or
								((vState = 80) and (hState = 594)) or
								((vState = 80) and (hState = 595)) or
								((vState = 81) and (hState = 455)) or
								((vState = 81) and (hState = 456)) or
								((vState = 81) and (hState = 457)) or
								((vState = 81) and (hState = 466)) or
								((vState = 81) and (hState = 467)) or
								((vState = 81) and (hState = 473)) or
								((vState = 81) and (hState = 474)) or
								((vState = 81) and (hState = 475)) or
								((vState = 81) and (hState = 476)) or
								((vState = 81) and (hState = 485)) or
								((vState = 81) and (hState = 486)) or
								((vState = 81) and (hState = 487)) or
								((vState = 81) and (hState = 488)) or
								((vState = 81) and (hState = 489)) or
								((vState = 81) and (hState = 490)) or
								((vState = 81) and (hState = 491)) or
								((vState = 81) and (hState = 492)) or
								((vState = 81) and (hState = 493)) or
								((vState = 81) and (hState = 494)) or
								((vState = 81) and (hState = 495)) or
								((vState = 81) and (hState = 496)) or
								((vState = 81) and (hState = 499)) or
								((vState = 81) and (hState = 500)) or
								((vState = 81) and (hState = 501)) or
								((vState = 81) and (hState = 504)) or
								((vState = 81) and (hState = 505)) or
								((vState = 81) and (hState = 507)) or
								((vState = 81) and (hState = 508)) or
								((vState = 81) and (hState = 509)) or
								((vState = 81) and (hState = 510)) or
								((vState = 81) and (hState = 511)) or
								((vState = 81) and (hState = 512)) or
								((vState = 81) and (hState = 513)) or
								((vState = 81) and (hState = 514)) or
								((vState = 81) and (hState = 515)) or
								((vState = 81) and (hState = 516)) or
								((vState = 81) and (hState = 517)) or
								((vState = 81) and (hState = 520)) or
								((vState = 81) and (hState = 523)) or
								((vState = 81) and (hState = 524)) or
								((vState = 81) and (hState = 525)) or
								((vState = 81) and (hState = 526)) or
								((vState = 81) and (hState = 527)) or
								((vState = 81) and (hState = 532)) or
								((vState = 81) and (hState = 533)) or
								((vState = 81) and (hState = 534)) or
								((vState = 81) and (hState = 544)) or
								((vState = 81) and (hState = 545)) or
								((vState = 81) and (hState = 546)) or
								((vState = 81) and (hState = 547)) or
								((vState = 81) and (hState = 548)) or
								((vState = 81) and (hState = 549)) or
								((vState = 81) and (hState = 550)) or
								((vState = 81) and (hState = 551)) or
								((vState = 81) and (hState = 552)) or
								((vState = 81) and (hState = 553)) or
								((vState = 81) and (hState = 554)) or
								((vState = 81) and (hState = 555)) or
								((vState = 81) and (hState = 556)) or
								((vState = 81) and (hState = 557)) or
								((vState = 81) and (hState = 558)) or
								((vState = 81) and (hState = 559)) or
								((vState = 81) and (hState = 560)) or
								((vState = 81) and (hState = 561)) or
								((vState = 81) and (hState = 565)) or
								((vState = 81) and (hState = 566)) or
								((vState = 81) and (hState = 567)) or
								((vState = 81) and (hState = 572)) or
								((vState = 81) and (hState = 573)) or
								((vState = 81) and (hState = 576)) or
								((vState = 81) and (hState = 577)) or
								((vState = 81) and (hState = 581)) or
								((vState = 81) and (hState = 582)) or
								((vState = 81) and (hState = 586)) or
								((vState = 81) and (hState = 587)) or
								((vState = 81) and (hState = 588)) or
								((vState = 81) and (hState = 589)) or
								((vState = 81) and (hState = 590)) or
								((vState = 81) and (hState = 591)) or
								((vState = 81) and (hState = 592)) or
								((vState = 81) and (hState = 593)) or
								((vState = 81) and (hState = 594)) or
								((vState = 81) and (hState = 595)) or
								((vState = 82) and (hState = 466)) or
								((vState = 82) and (hState = 467)) or
								((vState = 82) and (hState = 473)) or
								((vState = 82) and (hState = 474)) or
								((vState = 82) and (hState = 476)) or
								((vState = 82) and (hState = 477)) or
								((vState = 82) and (hState = 484)) or
								((vState = 82) and (hState = 485)) or
								((vState = 82) and (hState = 486)) or
								((vState = 82) and (hState = 487)) or
								((vState = 82) and (hState = 488)) or
								((vState = 82) and (hState = 489)) or
								((vState = 82) and (hState = 490)) or
								((vState = 82) and (hState = 493)) or
								((vState = 82) and (hState = 494)) or
								((vState = 82) and (hState = 495)) or
								((vState = 82) and (hState = 496)) or
								((vState = 82) and (hState = 500)) or
								((vState = 82) and (hState = 501)) or
								((vState = 82) and (hState = 502)) or
								((vState = 82) and (hState = 504)) or
								((vState = 82) and (hState = 505)) or
								((vState = 82) and (hState = 508)) or
								((vState = 82) and (hState = 509)) or
								((vState = 82) and (hState = 510)) or
								((vState = 82) and (hState = 511)) or
								((vState = 82) and (hState = 512)) or
								((vState = 82) and (hState = 513)) or
								((vState = 82) and (hState = 514)) or
								((vState = 82) and (hState = 515)) or
								((vState = 82) and (hState = 516)) or
								((vState = 82) and (hState = 520)) or
								((vState = 82) and (hState = 523)) or
								((vState = 82) and (hState = 524)) or
								((vState = 82) and (hState = 525)) or
								((vState = 82) and (hState = 526)) or
								((vState = 82) and (hState = 527)) or
								((vState = 82) and (hState = 532)) or
								((vState = 82) and (hState = 533)) or
								((vState = 82) and (hState = 534)) or
								((vState = 82) and (hState = 545)) or
								((vState = 82) and (hState = 546)) or
								((vState = 82) and (hState = 547)) or
								((vState = 82) and (hState = 548)) or
								((vState = 82) and (hState = 549)) or
								((vState = 82) and (hState = 550)) or
								((vState = 82) and (hState = 551)) or
								((vState = 82) and (hState = 552)) or
								((vState = 82) and (hState = 553)) or
								((vState = 82) and (hState = 554)) or
								((vState = 82) and (hState = 555)) or
								((vState = 82) and (hState = 556)) or
								((vState = 82) and (hState = 557)) or
								((vState = 82) and (hState = 558)) or
								((vState = 82) and (hState = 559)) or
								((vState = 82) and (hState = 560)) or
								((vState = 82) and (hState = 561)) or
								((vState = 82) and (hState = 562)) or
								((vState = 82) and (hState = 563)) or
								((vState = 82) and (hState = 564)) or
								((vState = 82) and (hState = 565)) or
								((vState = 82) and (hState = 566)) or
								((vState = 82) and (hState = 567)) or
								((vState = 82) and (hState = 568)) or
								((vState = 82) and (hState = 572)) or
								((vState = 82) and (hState = 573)) or
								((vState = 82) and (hState = 576)) or
								((vState = 82) and (hState = 577)) or
								((vState = 82) and (hState = 581)) or
								((vState = 82) and (hState = 582)) or
								((vState = 82) and (hState = 586)) or
								((vState = 82) and (hState = 587)) or
								((vState = 82) and (hState = 590)) or
								((vState = 82) and (hState = 591)) or
								((vState = 82) and (hState = 592)) or
								((vState = 82) and (hState = 593)) or
								((vState = 82) and (hState = 594)) or
								((vState = 82) and (hState = 595)) or
								((vState = 82) and (hState = 596)) or
								((vState = 82) and (hState = 597)) or
								((vState = 83) and (hState = 466)) or
								((vState = 83) and (hState = 467)) or
								((vState = 83) and (hState = 477)) or
								((vState = 83) and (hState = 478)) or
								((vState = 83) and (hState = 484)) or
								((vState = 83) and (hState = 485)) or
								((vState = 83) and (hState = 486)) or
								((vState = 83) and (hState = 494)) or
								((vState = 83) and (hState = 495)) or
								((vState = 83) and (hState = 496)) or
								((vState = 83) and (hState = 500)) or
								((vState = 83) and (hState = 501)) or
								((vState = 83) and (hState = 502)) or
								((vState = 83) and (hState = 504)) or
								((vState = 83) and (hState = 505)) or
								((vState = 83) and (hState = 509)) or
								((vState = 83) and (hState = 510)) or
								((vState = 83) and (hState = 511)) or
								((vState = 83) and (hState = 512)) or
								((vState = 83) and (hState = 513)) or
								((vState = 83) and (hState = 514)) or
								((vState = 83) and (hState = 515)) or
								((vState = 83) and (hState = 516)) or
								((vState = 83) and (hState = 520)) or
								((vState = 83) and (hState = 521)) or
								((vState = 83) and (hState = 522)) or
								((vState = 83) and (hState = 523)) or
								((vState = 83) and (hState = 524)) or
								((vState = 83) and (hState = 525)) or
								((vState = 83) and (hState = 526)) or
								((vState = 83) and (hState = 527)) or
								((vState = 83) and (hState = 528)) or
								((vState = 83) and (hState = 529)) or
								((vState = 83) and (hState = 530)) or
								((vState = 83) and (hState = 531)) or
								((vState = 83) and (hState = 532)) or
								((vState = 83) and (hState = 533)) or
								((vState = 83) and (hState = 534)) or
								((vState = 83) and (hState = 535)) or
								((vState = 83) and (hState = 536)) or
								((vState = 83) and (hState = 537)) or
								((vState = 83) and (hState = 538)) or
								((vState = 83) and (hState = 539)) or
								((vState = 83) and (hState = 546)) or
								((vState = 83) and (hState = 547)) or
								((vState = 83) and (hState = 548)) or
								((vState = 83) and (hState = 550)) or
								((vState = 83) and (hState = 551)) or
								((vState = 83) and (hState = 552)) or
								((vState = 83) and (hState = 553)) or
								((vState = 83) and (hState = 554)) or
								((vState = 83) and (hState = 555)) or
								((vState = 83) and (hState = 556)) or
								((vState = 83) and (hState = 557)) or
								((vState = 83) and (hState = 558)) or
								((vState = 83) and (hState = 559)) or
								((vState = 83) and (hState = 560)) or
								((vState = 83) and (hState = 561)) or
								((vState = 83) and (hState = 562)) or
								((vState = 83) and (hState = 563)) or
								((vState = 83) and (hState = 564)) or
								((vState = 83) and (hState = 566)) or
								((vState = 83) and (hState = 567)) or
								((vState = 83) and (hState = 568)) or
								((vState = 83) and (hState = 569)) or
								((vState = 83) and (hState = 572)) or
								((vState = 83) and (hState = 573)) or
								((vState = 83) and (hState = 575)) or
								((vState = 83) and (hState = 576)) or
								((vState = 83) and (hState = 577)) or
								((vState = 83) and (hState = 580)) or
								((vState = 83) and (hState = 581)) or
								((vState = 83) and (hState = 582)) or
								((vState = 83) and (hState = 586)) or
								((vState = 83) and (hState = 587)) or
								((vState = 83) and (hState = 591)) or
								((vState = 83) and (hState = 592)) or
								((vState = 83) and (hState = 593)) or
								((vState = 83) and (hState = 594)) or
								((vState = 83) and (hState = 596)) or
								((vState = 83) and (hState = 597)) or
								((vState = 83) and (hState = 598)) or
								((vState = 84) and (hState = 466)) or
								((vState = 84) and (hState = 467)) or
								((vState = 84) and (hState = 478)) or
								((vState = 84) and (hState = 479)) or
								((vState = 84) and (hState = 484)) or
								((vState = 84) and (hState = 485)) or
								((vState = 84) and (hState = 494)) or
								((vState = 84) and (hState = 495)) or
								((vState = 84) and (hState = 501)) or
								((vState = 84) and (hState = 502)) or
								((vState = 84) and (hState = 503)) or
								((vState = 84) and (hState = 504)) or
								((vState = 84) and (hState = 505)) or
								((vState = 84) and (hState = 510)) or
								((vState = 84) and (hState = 511)) or
								((vState = 84) and (hState = 512)) or
								((vState = 84) and (hState = 513)) or
								((vState = 84) and (hState = 514)) or
								((vState = 84) and (hState = 515)) or
								((vState = 84) and (hState = 516)) or
								((vState = 84) and (hState = 517)) or
								((vState = 84) and (hState = 520)) or
								((vState = 84) and (hState = 521)) or
								((vState = 84) and (hState = 522)) or
								((vState = 84) and (hState = 523)) or
								((vState = 84) and (hState = 527)) or
								((vState = 84) and (hState = 528)) or
								((vState = 84) and (hState = 531)) or
								((vState = 84) and (hState = 532)) or
								((vState = 84) and (hState = 533)) or
								((vState = 84) and (hState = 534)) or
								((vState = 84) and (hState = 535)) or
								((vState = 84) and (hState = 536)) or
								((vState = 84) and (hState = 537)) or
								((vState = 84) and (hState = 538)) or
								((vState = 84) and (hState = 539)) or
								((vState = 84) and (hState = 540)) or
								((vState = 84) and (hState = 541)) or
								((vState = 84) and (hState = 542)) or
								((vState = 84) and (hState = 543)) or
								((vState = 84) and (hState = 544)) or
								((vState = 84) and (hState = 545)) or
								((vState = 84) and (hState = 546)) or
								((vState = 84) and (hState = 547)) or
								((vState = 84) and (hState = 548)) or
								((vState = 84) and (hState = 549)) or
								((vState = 84) and (hState = 550)) or
								((vState = 84) and (hState = 551)) or
								((vState = 84) and (hState = 552)) or
								((vState = 84) and (hState = 553)) or
								((vState = 84) and (hState = 554)) or
								((vState = 84) and (hState = 555)) or
								((vState = 84) and (hState = 556)) or
								((vState = 84) and (hState = 557)) or
								((vState = 84) and (hState = 558)) or
								((vState = 84) and (hState = 559)) or
								((vState = 84) and (hState = 562)) or
								((vState = 84) and (hState = 563)) or
								((vState = 84) and (hState = 564)) or
								((vState = 84) and (hState = 567)) or
								((vState = 84) and (hState = 568)) or
								((vState = 84) and (hState = 569)) or
								((vState = 84) and (hState = 570)) or
								((vState = 84) and (hState = 572)) or
								((vState = 84) and (hState = 573)) or
								((vState = 84) and (hState = 574)) or
								((vState = 84) and (hState = 575)) or
								((vState = 84) and (hState = 576)) or
								((vState = 84) and (hState = 577)) or
								((vState = 84) and (hState = 580)) or
								((vState = 84) and (hState = 581)) or
								((vState = 84) and (hState = 582)) or
								((vState = 84) and (hState = 586)) or
								((vState = 84) and (hState = 587)) or
								((vState = 84) and (hState = 590)) or
								((vState = 84) and (hState = 591)) or
								((vState = 84) and (hState = 592)) or
								((vState = 84) and (hState = 593)) or
								((vState = 84) and (hState = 594)) or
								((vState = 84) and (hState = 597)) or
								((vState = 84) and (hState = 598)) or
								((vState = 84) and (hState = 599)) or
								((vState = 85) and (hState = 466)) or
								((vState = 85) and (hState = 467)) or
								((vState = 85) and (hState = 479)) or
								((vState = 85) and (hState = 480)) or
								((vState = 85) and (hState = 484)) or
								((vState = 85) and (hState = 485)) or
								((vState = 85) and (hState = 494)) or
								((vState = 85) and (hState = 495)) or
								((vState = 85) and (hState = 502)) or
								((vState = 85) and (hState = 503)) or
								((vState = 85) and (hState = 504)) or
								((vState = 85) and (hState = 505)) or
								((vState = 85) and (hState = 510)) or
								((vState = 85) and (hState = 511)) or
								((vState = 85) and (hState = 512)) or
								((vState = 85) and (hState = 513)) or
								((vState = 85) and (hState = 514)) or
								((vState = 85) and (hState = 515)) or
								((vState = 85) and (hState = 516)) or
								((vState = 85) and (hState = 517)) or
								((vState = 85) and (hState = 518)) or
								((vState = 85) and (hState = 519)) or
								((vState = 85) and (hState = 520)) or
								((vState = 85) and (hState = 521)) or
								((vState = 85) and (hState = 522)) or
								((vState = 85) and (hState = 523)) or
								((vState = 85) and (hState = 527)) or
								((vState = 85) and (hState = 528)) or
								((vState = 85) and (hState = 532)) or
								((vState = 85) and (hState = 533)) or
								((vState = 85) and (hState = 541)) or
								((vState = 85) and (hState = 542)) or
								((vState = 85) and (hState = 543)) or
								((vState = 85) and (hState = 544)) or
								((vState = 85) and (hState = 545)) or
								((vState = 85) and (hState = 546)) or
								((vState = 85) and (hState = 547)) or
								((vState = 85) and (hState = 548)) or
								((vState = 85) and (hState = 549)) or
								((vState = 85) and (hState = 550)) or
								((vState = 85) and (hState = 551)) or
								((vState = 85) and (hState = 552)) or
								((vState = 85) and (hState = 553)) or
								((vState = 85) and (hState = 554)) or
								((vState = 85) and (hState = 555)) or
								((vState = 85) and (hState = 556)) or
								((vState = 85) and (hState = 557)) or
								((vState = 85) and (hState = 563)) or
								((vState = 85) and (hState = 564)) or
								((vState = 85) and (hState = 565)) or
								((vState = 85) and (hState = 567)) or
								((vState = 85) and (hState = 568)) or
								((vState = 85) and (hState = 569)) or
								((vState = 85) and (hState = 570)) or
								((vState = 85) and (hState = 571)) or
								((vState = 85) and (hState = 572)) or
								((vState = 85) and (hState = 573)) or
								((vState = 85) and (hState = 574)) or
								((vState = 85) and (hState = 575)) or
								((vState = 85) and (hState = 576)) or
								((vState = 85) and (hState = 577)) or
								((vState = 85) and (hState = 580)) or
								((vState = 85) and (hState = 581)) or
								((vState = 85) and (hState = 582)) or
								((vState = 85) and (hState = 585)) or
								((vState = 85) and (hState = 586)) or
								((vState = 85) and (hState = 590)) or
								((vState = 85) and (hState = 591)) or
								((vState = 85) and (hState = 592)) or
								((vState = 85) and (hState = 593)) or
								((vState = 85) and (hState = 594)) or
								((vState = 85) and (hState = 598)) or
								((vState = 85) and (hState = 599)) or
								((vState = 86) and (hState = 467)) or
								((vState = 86) and (hState = 468)) or
								((vState = 86) and (hState = 479)) or
								((vState = 86) and (hState = 480)) or
								((vState = 86) and (hState = 481)) or
								((vState = 86) and (hState = 484)) or
								((vState = 86) and (hState = 485)) or
								((vState = 86) and (hState = 494)) or
								((vState = 86) and (hState = 495)) or
								((vState = 86) and (hState = 496)) or
								((vState = 86) and (hState = 503)) or
								((vState = 86) and (hState = 504)) or
								((vState = 86) and (hState = 505)) or
								((vState = 86) and (hState = 509)) or
								((vState = 86) and (hState = 510)) or
								((vState = 86) and (hState = 511)) or
								((vState = 86) and (hState = 512)) or
								((vState = 86) and (hState = 513)) or
								((vState = 86) and (hState = 514)) or
								((vState = 86) and (hState = 515)) or
								((vState = 86) and (hState = 518)) or
								((vState = 86) and (hState = 519)) or
								((vState = 86) and (hState = 520)) or
								((vState = 86) and (hState = 521)) or
								((vState = 86) and (hState = 522)) or
								((vState = 86) and (hState = 528)) or
								((vState = 86) and (hState = 531)) or
								((vState = 86) and (hState = 532)) or
								((vState = 86) and (hState = 544)) or
								((vState = 86) and (hState = 545)) or
								((vState = 86) and (hState = 546)) or
								((vState = 86) and (hState = 547)) or
								((vState = 86) and (hState = 548)) or
								((vState = 86) and (hState = 549)) or
								((vState = 86) and (hState = 550)) or
								((vState = 86) and (hState = 551)) or
								((vState = 86) and (hState = 552)) or
								((vState = 86) and (hState = 553)) or
								((vState = 86) and (hState = 554)) or
								((vState = 86) and (hState = 556)) or
								((vState = 86) and (hState = 557)) or
								((vState = 86) and (hState = 558)) or
								((vState = 86) and (hState = 559)) or
								((vState = 86) and (hState = 560)) or
								((vState = 86) and (hState = 561)) or
								((vState = 86) and (hState = 564)) or
								((vState = 86) and (hState = 565)) or
								((vState = 86) and (hState = 566)) or
								((vState = 86) and (hState = 567)) or
								((vState = 86) and (hState = 568)) or
								((vState = 86) and (hState = 569)) or
								((vState = 86) and (hState = 570)) or
								((vState = 86) and (hState = 571)) or
								((vState = 86) and (hState = 572)) or
								((vState = 86) and (hState = 573)) or
								((vState = 86) and (hState = 574)) or
								((vState = 86) and (hState = 575)) or
								((vState = 86) and (hState = 576)) or
								((vState = 86) and (hState = 577)) or
								((vState = 86) and (hState = 579)) or
								((vState = 86) and (hState = 580)) or
								((vState = 86) and (hState = 581)) or
								((vState = 86) and (hState = 585)) or
								((vState = 86) and (hState = 586)) or
								((vState = 86) and (hState = 589)) or
								((vState = 86) and (hState = 590)) or
								((vState = 86) and (hState = 592)) or
								((vState = 86) and (hState = 593)) or
								((vState = 86) and (hState = 594)) or
								((vState = 86) and (hState = 595)) or
								((vState = 86) and (hState = 599)) or
								((vState = 87) and (hState = 468)) or
								((vState = 87) and (hState = 469)) or
								((vState = 87) and (hState = 480)) or
								((vState = 87) and (hState = 481)) or
								((vState = 87) and (hState = 483)) or
								((vState = 87) and (hState = 484)) or
								((vState = 87) and (hState = 485)) or
								((vState = 87) and (hState = 494)) or
								((vState = 87) and (hState = 495)) or
								((vState = 87) and (hState = 496)) or
								((vState = 87) and (hState = 503)) or
								((vState = 87) and (hState = 504)) or
								((vState = 87) and (hState = 508)) or
								((vState = 87) and (hState = 509)) or
								((vState = 87) and (hState = 510)) or
								((vState = 87) and (hState = 511)) or
								((vState = 87) and (hState = 512)) or
								((vState = 87) and (hState = 513)) or
								((vState = 87) and (hState = 514)) or
								((vState = 87) and (hState = 515)) or
								((vState = 87) and (hState = 519)) or
								((vState = 87) and (hState = 520)) or
								((vState = 87) and (hState = 521)) or
								((vState = 87) and (hState = 522)) or
								((vState = 87) and (hState = 528)) or
								((vState = 87) and (hState = 529)) or
								((vState = 87) and (hState = 531)) or
								((vState = 87) and (hState = 532)) or
								((vState = 87) and (hState = 543)) or
								((vState = 87) and (hState = 544)) or
								((vState = 87) and (hState = 545)) or
								((vState = 87) and (hState = 546)) or
								((vState = 87) and (hState = 547)) or
								((vState = 87) and (hState = 548)) or
								((vState = 87) and (hState = 549)) or
								((vState = 87) and (hState = 550)) or
								((vState = 87) and (hState = 551)) or
								((vState = 87) and (hState = 552)) or
								((vState = 87) and (hState = 553)) or
								((vState = 87) and (hState = 554)) or
								((vState = 87) and (hState = 555)) or
								((vState = 87) and (hState = 556)) or
								((vState = 87) and (hState = 557)) or
								((vState = 87) and (hState = 558)) or
								((vState = 87) and (hState = 559)) or
								((vState = 87) and (hState = 560)) or
								((vState = 87) and (hState = 561)) or
								((vState = 87) and (hState = 562)) or
								((vState = 87) and (hState = 563)) or
								((vState = 87) and (hState = 564)) or
								((vState = 87) and (hState = 565)) or
								((vState = 87) and (hState = 566)) or
								((vState = 87) and (hState = 567)) or
								((vState = 87) and (hState = 568)) or
								((vState = 87) and (hState = 569)) or
								((vState = 87) and (hState = 570)) or
								((vState = 87) and (hState = 571)) or
								((vState = 87) and (hState = 572)) or
								((vState = 87) and (hState = 573)) or
								((vState = 87) and (hState = 574)) or
								((vState = 87) and (hState = 575)) or
								((vState = 87) and (hState = 576)) or
								((vState = 87) and (hState = 578)) or
								((vState = 87) and (hState = 579)) or
								((vState = 87) and (hState = 580)) or
								((vState = 87) and (hState = 581)) or
								((vState = 87) and (hState = 585)) or
								((vState = 87) and (hState = 586)) or
								((vState = 87) and (hState = 588)) or
								((vState = 87) and (hState = 589)) or
								((vState = 87) and (hState = 593)) or
								((vState = 87) and (hState = 594)) or
								((vState = 87) and (hState = 595)) or
								((vState = 87) and (hState = 596)) or
								((vState = 88) and (hState = 468)) or
								((vState = 88) and (hState = 469)) or
								((vState = 88) and (hState = 481)) or
								((vState = 88) and (hState = 482)) or
								((vState = 88) and (hState = 483)) or
								((vState = 88) and (hState = 484)) or
								((vState = 88) and (hState = 485)) or
								((vState = 88) and (hState = 489)) or
								((vState = 88) and (hState = 494)) or
								((vState = 88) and (hState = 495)) or
								((vState = 88) and (hState = 496)) or
								((vState = 88) and (hState = 497)) or
								((vState = 88) and (hState = 503)) or
								((vState = 88) and (hState = 504)) or
								((vState = 88) and (hState = 508)) or
								((vState = 88) and (hState = 509)) or
								((vState = 88) and (hState = 510)) or
								((vState = 88) and (hState = 511)) or
								((vState = 88) and (hState = 512)) or
								((vState = 88) and (hState = 514)) or
								((vState = 88) and (hState = 515)) or
								((vState = 88) and (hState = 516)) or
								((vState = 88) and (hState = 520)) or
								((vState = 88) and (hState = 521)) or
								((vState = 88) and (hState = 522)) or
								((vState = 88) and (hState = 528)) or
								((vState = 88) and (hState = 529)) or
								((vState = 88) and (hState = 531)) or
								((vState = 88) and (hState = 532)) or
								((vState = 88) and (hState = 542)) or
								((vState = 88) and (hState = 543)) or
								((vState = 88) and (hState = 544)) or
								((vState = 88) and (hState = 545)) or
								((vState = 88) and (hState = 546)) or
								((vState = 88) and (hState = 547)) or
								((vState = 88) and (hState = 548)) or
								((vState = 88) and (hState = 549)) or
								((vState = 88) and (hState = 550)) or
								((vState = 88) and (hState = 551)) or
								((vState = 88) and (hState = 554)) or
								((vState = 88) and (hState = 555)) or
								((vState = 88) and (hState = 556)) or
								((vState = 88) and (hState = 558)) or
								((vState = 88) and (hState = 559)) or
								((vState = 88) and (hState = 563)) or
								((vState = 88) and (hState = 564)) or
								((vState = 88) and (hState = 565)) or
								((vState = 88) and (hState = 566)) or
								((vState = 88) and (hState = 567)) or
								((vState = 88) and (hState = 568)) or
								((vState = 88) and (hState = 569)) or
								((vState = 88) and (hState = 570)) or
								((vState = 88) and (hState = 571)) or
								((vState = 88) and (hState = 572)) or
								((vState = 88) and (hState = 573)) or
								((vState = 88) and (hState = 574)) or
								((vState = 88) and (hState = 575)) or
								((vState = 88) and (hState = 576)) or
								((vState = 88) and (hState = 577)) or
								((vState = 88) and (hState = 578)) or
								((vState = 88) and (hState = 579)) or
								((vState = 88) and (hState = 580)) or
								((vState = 88) and (hState = 581)) or
								((vState = 88) and (hState = 584)) or
								((vState = 88) and (hState = 585)) or
								((vState = 88) and (hState = 586)) or
								((vState = 88) and (hState = 587)) or
								((vState = 88) and (hState = 588)) or
								((vState = 88) and (hState = 593)) or
								((vState = 88) and (hState = 594)) or
								((vState = 88) and (hState = 595)) or
								((vState = 88) and (hState = 596)) or
								((vState = 88) and (hState = 597)) or
								((vState = 88) and (hState = 599)) or
								((vState = 89) and (hState = 469)) or
								((vState = 89) and (hState = 470)) or
								((vState = 89) and (hState = 481)) or
								((vState = 89) and (hState = 482)) or
								((vState = 89) and (hState = 483)) or
								((vState = 89) and (hState = 484)) or
								((vState = 89) and (hState = 485)) or
								((vState = 89) and (hState = 489)) or
								((vState = 89) and (hState = 490)) or
								((vState = 89) and (hState = 493)) or
								((vState = 89) and (hState = 494)) or
								((vState = 89) and (hState = 495)) or
								((vState = 89) and (hState = 496)) or
								((vState = 89) and (hState = 497)) or
								((vState = 89) and (hState = 503)) or
								((vState = 89) and (hState = 508)) or
								((vState = 89) and (hState = 509)) or
								((vState = 89) and (hState = 510)) or
								((vState = 89) and (hState = 511)) or
								((vState = 89) and (hState = 515)) or
								((vState = 89) and (hState = 516)) or
								((vState = 89) and (hState = 517)) or
								((vState = 89) and (hState = 521)) or
								((vState = 89) and (hState = 529)) or
								((vState = 89) and (hState = 530)) or
								((vState = 89) and (hState = 531)) or
								((vState = 89) and (hState = 532)) or
								((vState = 89) and (hState = 537)) or
								((vState = 89) and (hState = 538)) or
								((vState = 89) and (hState = 539)) or
								((vState = 89) and (hState = 540)) or
								((vState = 89) and (hState = 541)) or
								((vState = 89) and (hState = 542)) or
								((vState = 89) and (hState = 543)) or
								((vState = 89) and (hState = 544)) or
								((vState = 89) and (hState = 545)) or
								((vState = 89) and (hState = 546)) or
								((vState = 89) and (hState = 547)) or
								((vState = 89) and (hState = 548)) or
								((vState = 89) and (hState = 549)) or
								((vState = 89) and (hState = 555)) or
								((vState = 89) and (hState = 556)) or
								((vState = 89) and (hState = 559)) or
								((vState = 89) and (hState = 560)) or
								((vState = 89) and (hState = 564)) or
								((vState = 89) and (hState = 565)) or
								((vState = 89) and (hState = 566)) or
								((vState = 89) and (hState = 567)) or
								((vState = 89) and (hState = 568)) or
								((vState = 89) and (hState = 569)) or
								((vState = 89) and (hState = 570)) or
								((vState = 89) and (hState = 571)) or
								((vState = 89) and (hState = 572)) or
								((vState = 89) and (hState = 573)) or
								((vState = 89) and (hState = 575)) or
								((vState = 89) and (hState = 576)) or
								((vState = 89) and (hState = 577)) or
								((vState = 89) and (hState = 578)) or
								((vState = 89) and (hState = 579)) or
								((vState = 89) and (hState = 580)) or
								((vState = 89) and (hState = 581)) or
								((vState = 89) and (hState = 584)) or
								((vState = 89) and (hState = 585)) or
								((vState = 89) and (hState = 586)) or
								((vState = 89) and (hState = 587)) or
								((vState = 89) and (hState = 588)) or
								((vState = 89) and (hState = 593)) or
								((vState = 89) and (hState = 594)) or
								((vState = 89) and (hState = 595)) or
								((vState = 89) and (hState = 596)) or
								((vState = 89) and (hState = 597)) or
								((vState = 89) and (hState = 598)) or
								((vState = 89) and (hState = 599)) or
								((vState = 90) and (hState = 469)) or
								((vState = 90) and (hState = 470)) or
								((vState = 90) and (hState = 482)) or
								((vState = 90) and (hState = 483)) or
								((vState = 90) and (hState = 484)) or
								((vState = 90) and (hState = 485)) or
								((vState = 90) and (hState = 489)) or
								((vState = 90) and (hState = 490)) or
								((vState = 90) and (hState = 491)) or
								((vState = 90) and (hState = 493)) or
								((vState = 90) and (hState = 494)) or
								((vState = 90) and (hState = 496)) or
								((vState = 90) and (hState = 497)) or
								((vState = 90) and (hState = 500)) or
								((vState = 90) and (hState = 501)) or
								((vState = 90) and (hState = 502)) or
								((vState = 90) and (hState = 503)) or
								((vState = 90) and (hState = 509)) or
								((vState = 90) and (hState = 510)) or
								((vState = 90) and (hState = 511)) or
								((vState = 90) and (hState = 515)) or
								((vState = 90) and (hState = 516)) or
								((vState = 90) and (hState = 517)) or
								((vState = 90) and (hState = 518)) or
								((vState = 90) and (hState = 521)) or
								((vState = 90) and (hState = 522)) or
								((vState = 90) and (hState = 529)) or
								((vState = 90) and (hState = 530)) or
								((vState = 90) and (hState = 531)) or
								((vState = 90) and (hState = 537)) or
								((vState = 90) and (hState = 538)) or
								((vState = 90) and (hState = 539)) or
								((vState = 90) and (hState = 540)) or
								((vState = 90) and (hState = 541)) or
								((vState = 90) and (hState = 542)) or
								((vState = 90) and (hState = 549)) or
								((vState = 90) and (hState = 554)) or
								((vState = 90) and (hState = 555)) or
								((vState = 90) and (hState = 556)) or
								((vState = 90) and (hState = 557)) or
								((vState = 90) and (hState = 559)) or
								((vState = 90) and (hState = 560)) or
								((vState = 90) and (hState = 563)) or
								((vState = 90) and (hState = 564)) or
								((vState = 90) and (hState = 565)) or
								((vState = 90) and (hState = 566)) or
								((vState = 90) and (hState = 567)) or
								((vState = 90) and (hState = 568)) or
								((vState = 90) and (hState = 569)) or
								((vState = 90) and (hState = 570)) or
								((vState = 90) and (hState = 571)) or
								((vState = 90) and (hState = 572)) or
								((vState = 90) and (hState = 573)) or
								((vState = 90) and (hState = 575)) or
								((vState = 90) and (hState = 576)) or
								((vState = 90) and (hState = 577)) or
								((vState = 90) and (hState = 579)) or
								((vState = 90) and (hState = 580)) or
								((vState = 90) and (hState = 581)) or
								((vState = 90) and (hState = 584)) or
								((vState = 90) and (hState = 585)) or
								((vState = 90) and (hState = 586)) or
								((vState = 90) and (hState = 587)) or
								((vState = 90) and (hState = 593)) or
								((vState = 90) and (hState = 594)) or
								((vState = 90) and (hState = 595)) or
								((vState = 90) and (hState = 598)) or
								((vState = 90) and (hState = 599)) or
								((vState = 91) and (hState = 470)) or
								((vState = 91) and (hState = 471)) or
								((vState = 91) and (hState = 477)) or
								((vState = 91) and (hState = 482)) or
								((vState = 91) and (hState = 483)) or
								((vState = 91) and (hState = 484)) or
								((vState = 91) and (hState = 485)) or
								((vState = 91) and (hState = 488)) or
								((vState = 91) and (hState = 489)) or
								((vState = 91) and (hState = 490)) or
								((vState = 91) and (hState = 491)) or
								((vState = 91) and (hState = 493)) or
								((vState = 91) and (hState = 494)) or
								((vState = 91) and (hState = 496)) or
								((vState = 91) and (hState = 497)) or
								((vState = 91) and (hState = 498)) or
								((vState = 91) and (hState = 499)) or
								((vState = 91) and (hState = 500)) or
								((vState = 91) and (hState = 501)) or
								((vState = 91) and (hState = 502)) or
								((vState = 91) and (hState = 503)) or
								((vState = 91) and (hState = 508)) or
								((vState = 91) and (hState = 509)) or
								((vState = 91) and (hState = 510)) or
								((vState = 91) and (hState = 511)) or
								((vState = 91) and (hState = 512)) or
								((vState = 91) and (hState = 513)) or
								((vState = 91) and (hState = 515)) or
								((vState = 91) and (hState = 516)) or
								((vState = 91) and (hState = 517)) or
								((vState = 91) and (hState = 518)) or
								((vState = 91) and (hState = 519)) or
								((vState = 91) and (hState = 521)) or
								((vState = 91) and (hState = 522)) or
								((vState = 91) and (hState = 529)) or
								((vState = 91) and (hState = 530)) or
								((vState = 91) and (hState = 531)) or
								((vState = 91) and (hState = 536)) or
								((vState = 91) and (hState = 537)) or
								((vState = 91) and (hState = 538)) or
								((vState = 91) and (hState = 539)) or
								((vState = 91) and (hState = 540)) or
								((vState = 91) and (hState = 541)) or
								((vState = 91) and (hState = 542)) or
								((vState = 91) and (hState = 543)) or
								((vState = 91) and (hState = 544)) or
								((vState = 91) and (hState = 549)) or
								((vState = 91) and (hState = 554)) or
								((vState = 91) and (hState = 555)) or
								((vState = 91) and (hState = 556)) or
								((vState = 91) and (hState = 557)) or
								((vState = 91) and (hState = 558)) or
								((vState = 91) and (hState = 560)) or
								((vState = 91) and (hState = 561)) or
								((vState = 91) and (hState = 562)) or
								((vState = 91) and (hState = 563)) or
								((vState = 91) and (hState = 564)) or
								((vState = 91) and (hState = 565)) or
								((vState = 91) and (hState = 566)) or
								((vState = 91) and (hState = 567)) or
								((vState = 91) and (hState = 568)) or
								((vState = 91) and (hState = 569)) or
								((vState = 91) and (hState = 570)) or
								((vState = 91) and (hState = 571)) or
								((vState = 91) and (hState = 572)) or
								((vState = 91) and (hState = 573)) or
								((vState = 91) and (hState = 574)) or
								((vState = 91) and (hState = 575)) or
								((vState = 91) and (hState = 576)) or
								((vState = 91) and (hState = 578)) or
								((vState = 91) and (hState = 579)) or
								((vState = 91) and (hState = 580)) or
								((vState = 91) and (hState = 581)) or
								((vState = 91) and (hState = 583)) or
								((vState = 91) and (hState = 584)) or
								((vState = 91) and (hState = 585)) or
								((vState = 91) and (hState = 586)) or
								((vState = 91) and (hState = 593)) or
								((vState = 91) and (hState = 594)) or
								((vState = 91) and (hState = 595)) or
								((vState = 91) and (hState = 596)) or
								((vState = 91) and (hState = 598)) or
								((vState = 91) and (hState = 599)) or
								((vState = 92) and (hState = 470)) or
								((vState = 92) and (hState = 471)) or
								((vState = 92) and (hState = 475)) or
								((vState = 92) and (hState = 476)) or
								((vState = 92) and (hState = 477)) or
								((vState = 92) and (hState = 478)) or
								((vState = 92) and (hState = 481)) or
								((vState = 92) and (hState = 482)) or
								((vState = 92) and (hState = 483)) or
								((vState = 92) and (hState = 484)) or
								((vState = 92) and (hState = 485)) or
								((vState = 92) and (hState = 488)) or
								((vState = 92) and (hState = 489)) or
								((vState = 92) and (hState = 491)) or
								((vState = 92) and (hState = 492)) or
								((vState = 92) and (hState = 493)) or
								((vState = 92) and (hState = 494)) or
								((vState = 92) and (hState = 495)) or
								((vState = 92) and (hState = 496)) or
								((vState = 92) and (hState = 497)) or
								((vState = 92) and (hState = 498)) or
								((vState = 92) and (hState = 499)) or
								((vState = 92) and (hState = 501)) or
								((vState = 92) and (hState = 502)) or
								((vState = 92) and (hState = 503)) or
								((vState = 92) and (hState = 508)) or
								((vState = 92) and (hState = 509)) or
								((vState = 92) and (hState = 512)) or
								((vState = 92) and (hState = 513)) or
								((vState = 92) and (hState = 514)) or
								((vState = 92) and (hState = 515)) or
								((vState = 92) and (hState = 516)) or
								((vState = 92) and (hState = 518)) or
								((vState = 92) and (hState = 519)) or
								((vState = 92) and (hState = 520)) or
								((vState = 92) and (hState = 521)) or
								((vState = 92) and (hState = 522)) or
								((vState = 92) and (hState = 529)) or
								((vState = 92) and (hState = 530)) or
								((vState = 92) and (hState = 531)) or
								((vState = 92) and (hState = 532)) or
								((vState = 92) and (hState = 533)) or
								((vState = 92) and (hState = 534)) or
								((vState = 92) and (hState = 535)) or
								((vState = 92) and (hState = 536)) or
								((vState = 92) and (hState = 537)) or
								((vState = 92) and (hState = 538)) or
								((vState = 92) and (hState = 539)) or
								((vState = 92) and (hState = 540)) or
								((vState = 92) and (hState = 541)) or
								((vState = 92) and (hState = 542)) or
								((vState = 92) and (hState = 543)) or
								((vState = 92) and (hState = 544)) or
								((vState = 92) and (hState = 545)) or
								((vState = 92) and (hState = 548)) or
								((vState = 92) and (hState = 549)) or
								((vState = 92) and (hState = 554)) or
								((vState = 92) and (hState = 555)) or
								((vState = 92) and (hState = 557)) or
								((vState = 92) and (hState = 558)) or
								((vState = 92) and (hState = 559)) or
								((vState = 92) and (hState = 560)) or
								((vState = 92) and (hState = 561)) or
								((vState = 92) and (hState = 562)) or
								((vState = 92) and (hState = 563)) or
								((vState = 92) and (hState = 564)) or
								((vState = 92) and (hState = 565)) or
								((vState = 92) and (hState = 566)) or
								((vState = 92) and (hState = 568)) or
								((vState = 92) and (hState = 569)) or
								((vState = 92) and (hState = 570)) or
								((vState = 92) and (hState = 571)) or
								((vState = 92) and (hState = 572)) or
								((vState = 92) and (hState = 573)) or
								((vState = 92) and (hState = 574)) or
								((vState = 92) and (hState = 575)) or
								((vState = 92) and (hState = 576)) or
								((vState = 92) and (hState = 578)) or
								((vState = 92) and (hState = 579)) or
								((vState = 92) and (hState = 580)) or
								((vState = 92) and (hState = 583)) or
								((vState = 92) and (hState = 584)) or
								((vState = 92) and (hState = 585)) or
								((vState = 92) and (hState = 586)) or
								((vState = 92) and (hState = 594)) or
								((vState = 92) and (hState = 595)) or
								((vState = 92) and (hState = 596)) or
								((vState = 92) and (hState = 598)) or
								((vState = 92) and (hState = 599)) or
								((vState = 93) and (hState = 471)) or
								((vState = 93) and (hState = 472)) or
								((vState = 93) and (hState = 474)) or
								((vState = 93) and (hState = 475)) or
								((vState = 93) and (hState = 476)) or
								((vState = 93) and (hState = 477)) or
								((vState = 93) and (hState = 478)) or
								((vState = 93) and (hState = 480)) or
								((vState = 93) and (hState = 481)) or
								((vState = 93) and (hState = 482)) or
								((vState = 93) and (hState = 483)) or
								((vState = 93) and (hState = 484)) or
								((vState = 93) and (hState = 485)) or
								((vState = 93) and (hState = 486)) or
								((vState = 93) and (hState = 488)) or
								((vState = 93) and (hState = 489)) or
								((vState = 93) and (hState = 491)) or
								((vState = 93) and (hState = 492)) or
								((vState = 93) and (hState = 493)) or
								((vState = 93) and (hState = 494)) or
								((vState = 93) and (hState = 495)) or
								((vState = 93) and (hState = 496)) or
								((vState = 93) and (hState = 498)) or
								((vState = 93) and (hState = 499)) or
								((vState = 93) and (hState = 501)) or
								((vState = 93) and (hState = 502)) or
								((vState = 93) and (hState = 503)) or
								((vState = 93) and (hState = 507)) or
								((vState = 93) and (hState = 508)) or
								((vState = 93) and (hState = 513)) or
								((vState = 93) and (hState = 514)) or
								((vState = 93) and (hState = 515)) or
								((vState = 93) and (hState = 516)) or
								((vState = 93) and (hState = 517)) or
								((vState = 93) and (hState = 519)) or
								((vState = 93) and (hState = 520)) or
								((vState = 93) and (hState = 521)) or
								((vState = 93) and (hState = 522)) or
								((vState = 93) and (hState = 523)) or
								((vState = 93) and (hState = 524)) or
								((vState = 93) and (hState = 526)) or
								((vState = 93) and (hState = 527)) or
								((vState = 93) and (hState = 528)) or
								((vState = 93) and (hState = 529)) or
								((vState = 93) and (hState = 530)) or
								((vState = 93) and (hState = 531)) or
								((vState = 93) and (hState = 532)) or
								((vState = 93) and (hState = 533)) or
								((vState = 93) and (hState = 534)) or
								((vState = 93) and (hState = 535)) or
								((vState = 93) and (hState = 536)) or
								((vState = 93) and (hState = 537)) or
								((vState = 93) and (hState = 538)) or
								((vState = 93) and (hState = 539)) or
								((vState = 93) and (hState = 540)) or
								((vState = 93) and (hState = 544)) or
								((vState = 93) and (hState = 545)) or
								((vState = 93) and (hState = 548)) or
								((vState = 93) and (hState = 549)) or
								((vState = 93) and (hState = 554)) or
								((vState = 93) and (hState = 555)) or
								((vState = 93) and (hState = 558)) or
								((vState = 93) and (hState = 559)) or
								((vState = 93) and (hState = 560)) or
								((vState = 93) and (hState = 561)) or
								((vState = 93) and (hState = 562)) or
								((vState = 93) and (hState = 563)) or
								((vState = 93) and (hState = 564)) or
								((vState = 93) and (hState = 565)) or
								((vState = 93) and (hState = 568)) or
								((vState = 93) and (hState = 569)) or
								((vState = 93) and (hState = 570)) or
								((vState = 93) and (hState = 571)) or
								((vState = 93) and (hState = 572)) or
								((vState = 93) and (hState = 573)) or
								((vState = 93) and (hState = 574)) or
								((vState = 93) and (hState = 575)) or
								((vState = 93) and (hState = 576)) or
								((vState = 93) and (hState = 578)) or
								((vState = 93) and (hState = 579)) or
								((vState = 93) and (hState = 580)) or
								((vState = 93) and (hState = 582)) or
								((vState = 93) and (hState = 583)) or
								((vState = 93) and (hState = 584)) or
								((vState = 93) and (hState = 586)) or
								((vState = 93) and (hState = 587)) or
								((vState = 93) and (hState = 594)) or
								((vState = 93) and (hState = 595)) or
								((vState = 93) and (hState = 596)) or
								((vState = 93) and (hState = 598)) or
								((vState = 93) and (hState = 599)) or
								((vState = 94) and (hState = 471)) or
								((vState = 94) and (hState = 472)) or
								((vState = 94) and (hState = 473)) or
								((vState = 94) and (hState = 474)) or
								((vState = 94) and (hState = 475)) or
								((vState = 94) and (hState = 477)) or
								((vState = 94) and (hState = 478)) or
								((vState = 94) and (hState = 480)) or
								((vState = 94) and (hState = 481)) or
								((vState = 94) and (hState = 482)) or
								((vState = 94) and (hState = 483)) or
								((vState = 94) and (hState = 484)) or
								((vState = 94) and (hState = 485)) or
								((vState = 94) and (hState = 486)) or
								((vState = 94) and (hState = 487)) or
								((vState = 94) and (hState = 488)) or
								((vState = 94) and (hState = 492)) or
								((vState = 94) and (hState = 493)) or
								((vState = 94) and (hState = 498)) or
								((vState = 94) and (hState = 499)) or
								((vState = 94) and (hState = 501)) or
								((vState = 94) and (hState = 502)) or
								((vState = 94) and (hState = 503)) or
								((vState = 94) and (hState = 505)) or
								((vState = 94) and (hState = 506)) or
								((vState = 94) and (hState = 507)) or
								((vState = 94) and (hState = 513)) or
								((vState = 94) and (hState = 514)) or
								((vState = 94) and (hState = 515)) or
								((vState = 94) and (hState = 516)) or
								((vState = 94) and (hState = 517)) or
								((vState = 94) and (hState = 518)) or
								((vState = 94) and (hState = 521)) or
								((vState = 94) and (hState = 522)) or
								((vState = 94) and (hState = 523)) or
								((vState = 94) and (hState = 524)) or
								((vState = 94) and (hState = 525)) or
								((vState = 94) and (hState = 526)) or
								((vState = 94) and (hState = 527)) or
								((vState = 94) and (hState = 528)) or
								((vState = 94) and (hState = 529)) or
								((vState = 94) and (hState = 530)) or
								((vState = 94) and (hState = 531)) or
								((vState = 94) and (hState = 532)) or
								((vState = 94) and (hState = 533)) or
								((vState = 94) and (hState = 534)) or
								((vState = 94) and (hState = 535)) or
								((vState = 94) and (hState = 536)) or
								((vState = 94) and (hState = 537)) or
								((vState = 94) and (hState = 538)) or
								((vState = 94) and (hState = 539)) or
								((vState = 94) and (hState = 545)) or
								((vState = 94) and (hState = 546)) or
								((vState = 94) and (hState = 548)) or
								((vState = 94) and (hState = 549)) or
								((vState = 94) and (hState = 555)) or
								((vState = 94) and (hState = 556)) or
								((vState = 94) and (hState = 557)) or
								((vState = 94) and (hState = 558)) or
								((vState = 94) and (hState = 559)) or
								((vState = 94) and (hState = 560)) or
								((vState = 94) and (hState = 561)) or
								((vState = 94) and (hState = 562)) or
								((vState = 94) and (hState = 563)) or
								((vState = 94) and (hState = 569)) or
								((vState = 94) and (hState = 570)) or
								((vState = 94) and (hState = 571)) or
								((vState = 94) and (hState = 572)) or
								((vState = 94) and (hState = 574)) or
								((vState = 94) and (hState = 575)) or
								((vState = 94) and (hState = 576)) or
								((vState = 94) and (hState = 577)) or
								((vState = 94) and (hState = 578)) or
								((vState = 94) and (hState = 579)) or
								((vState = 94) and (hState = 582)) or
								((vState = 94) and (hState = 583)) or
								((vState = 94) and (hState = 584)) or
								((vState = 94) and (hState = 586)) or
								((vState = 94) and (hState = 587)) or
								((vState = 94) and (hState = 593)) or
								((vState = 94) and (hState = 594)) or
								((vState = 94) and (hState = 595)) or
								((vState = 94) and (hState = 596)) or
								((vState = 94) and (hState = 598)) or
								((vState = 94) and (hState = 599)) or
								((vState = 95) and (hState = 472)) or
								((vState = 95) and (hState = 473)) or
								((vState = 95) and (hState = 474)) or
								((vState = 95) and (hState = 477)) or
								((vState = 95) and (hState = 478)) or
								((vState = 95) and (hState = 479)) or
								((vState = 95) and (hState = 480)) or
								((vState = 95) and (hState = 481)) or
								((vState = 95) and (hState = 482)) or
								((vState = 95) and (hState = 483)) or
								((vState = 95) and (hState = 484)) or
								((vState = 95) and (hState = 485)) or
								((vState = 95) and (hState = 486)) or
								((vState = 95) and (hState = 487)) or
								((vState = 95) and (hState = 488)) or
								((vState = 95) and (hState = 493)) or
								((vState = 95) and (hState = 494)) or
								((vState = 95) and (hState = 498)) or
								((vState = 95) and (hState = 499)) or
								((vState = 95) and (hState = 500)) or
								((vState = 95) and (hState = 501)) or
								((vState = 95) and (hState = 502)) or
								((vState = 95) and (hState = 503)) or
								((vState = 95) and (hState = 504)) or
								((vState = 95) and (hState = 505)) or
								((vState = 95) and (hState = 506)) or
								((vState = 95) and (hState = 512)) or
								((vState = 95) and (hState = 513)) or
								((vState = 95) and (hState = 516)) or
								((vState = 95) and (hState = 517)) or
								((vState = 95) and (hState = 518)) or
								((vState = 95) and (hState = 521)) or
								((vState = 95) and (hState = 522)) or
								((vState = 95) and (hState = 527)) or
								((vState = 95) and (hState = 528)) or
								((vState = 95) and (hState = 529)) or
								((vState = 95) and (hState = 530)) or
								((vState = 95) and (hState = 531)) or
								((vState = 95) and (hState = 532)) or
								((vState = 95) and (hState = 533)) or
								((vState = 95) and (hState = 534)) or
								((vState = 95) and (hState = 535)) or
								((vState = 95) and (hState = 536)) or
								((vState = 95) and (hState = 537)) or
								((vState = 95) and (hState = 538)) or
								((vState = 95) and (hState = 546)) or
								((vState = 95) and (hState = 547)) or
								((vState = 95) and (hState = 548)) or
								((vState = 95) and (hState = 555)) or
								((vState = 95) and (hState = 556)) or
								((vState = 95) and (hState = 557)) or
								((vState = 95) and (hState = 559)) or
								((vState = 95) and (hState = 560)) or
								((vState = 95) and (hState = 561)) or
								((vState = 95) and (hState = 562)) or
								((vState = 95) and (hState = 563)) or
								((vState = 95) and (hState = 564)) or
								((vState = 95) and (hState = 569)) or
								((vState = 95) and (hState = 570)) or
								((vState = 95) and (hState = 571)) or
								((vState = 95) and (hState = 572)) or
								((vState = 95) and (hState = 574)) or
								((vState = 95) and (hState = 575)) or
								((vState = 95) and (hState = 576)) or
								((vState = 95) and (hState = 577)) or
								((vState = 95) and (hState = 578)) or
								((vState = 95) and (hState = 579)) or
								((vState = 95) and (hState = 582)) or
								((vState = 95) and (hState = 583)) or
								((vState = 95) and (hState = 584)) or
								((vState = 95) and (hState = 586)) or
								((vState = 95) and (hState = 587)) or
								((vState = 95) and (hState = 593)) or
								((vState = 95) and (hState = 594)) or
								((vState = 95) and (hState = 596)) or
								((vState = 95) and (hState = 597)) or
								((vState = 95) and (hState = 598)) or
								((vState = 95) and (hState = 599)) or
								((vState = 96) and (hState = 470)) or
								((vState = 96) and (hState = 471)) or
								((vState = 96) and (hState = 472)) or
								((vState = 96) and (hState = 473)) or
								((vState = 96) and (hState = 474)) or
								((vState = 96) and (hState = 477)) or
								((vState = 96) and (hState = 478)) or
								((vState = 96) and (hState = 479)) or
								((vState = 96) and (hState = 480)) or
								((vState = 96) and (hState = 481)) or
								((vState = 96) and (hState = 482)) or
								((vState = 96) and (hState = 483)) or
								((vState = 96) and (hState = 484)) or
								((vState = 96) and (hState = 485)) or
								((vState = 96) and (hState = 486)) or
								((vState = 96) and (hState = 487)) or
								((vState = 96) and (hState = 488)) or
								((vState = 96) and (hState = 493)) or
								((vState = 96) and (hState = 494)) or
								((vState = 96) and (hState = 499)) or
								((vState = 96) and (hState = 500)) or
								((vState = 96) and (hState = 502)) or
								((vState = 96) and (hState = 503)) or
								((vState = 96) and (hState = 504)) or
								((vState = 96) and (hState = 505)) or
								((vState = 96) and (hState = 510)) or
								((vState = 96) and (hState = 511)) or
								((vState = 96) and (hState = 512)) or
								((vState = 96) and (hState = 516)) or
								((vState = 96) and (hState = 517)) or
								((vState = 96) and (hState = 518)) or
								((vState = 96) and (hState = 519)) or
								((vState = 96) and (hState = 520)) or
								((vState = 96) and (hState = 521)) or
								((vState = 96) and (hState = 522)) or
								((vState = 96) and (hState = 527)) or
								((vState = 96) and (hState = 528)) or
								((vState = 96) and (hState = 529)) or
								((vState = 96) and (hState = 533)) or
								((vState = 96) and (hState = 534)) or
								((vState = 96) and (hState = 535)) or
								((vState = 96) and (hState = 536)) or
								((vState = 96) and (hState = 537)) or
								((vState = 96) and (hState = 538)) or
								((vState = 96) and (hState = 539)) or
								((vState = 96) and (hState = 540)) or
								((vState = 96) and (hState = 541)) or
								((vState = 96) and (hState = 542)) or
								((vState = 96) and (hState = 543)) or
								((vState = 96) and (hState = 546)) or
								((vState = 96) and (hState = 547)) or
								((vState = 96) and (hState = 548)) or
								((vState = 96) and (hState = 554)) or
								((vState = 96) and (hState = 555)) or
								((vState = 96) and (hState = 556)) or
								((vState = 96) and (hState = 557)) or
								((vState = 96) and (hState = 558)) or
								((vState = 96) and (hState = 559)) or
								((vState = 96) and (hState = 560)) or
								((vState = 96) and (hState = 561)) or
								((vState = 96) and (hState = 562)) or
								((vState = 96) and (hState = 563)) or
								((vState = 96) and (hState = 564)) or
								((vState = 96) and (hState = 565)) or
								((vState = 96) and (hState = 568)) or
								((vState = 96) and (hState = 569)) or
								((vState = 96) and (hState = 570)) or
								((vState = 96) and (hState = 571)) or
								((vState = 96) and (hState = 572)) or
								((vState = 96) and (hState = 573)) or
								((vState = 96) and (hState = 574)) or
								((vState = 96) and (hState = 575)) or
								((vState = 96) and (hState = 576)) or
								((vState = 96) and (hState = 577)) or
								((vState = 96) and (hState = 578)) or
								((vState = 96) and (hState = 579)) or
								((vState = 96) and (hState = 581)) or
								((vState = 96) and (hState = 582)) or
								((vState = 96) and (hState = 583)) or
								((vState = 96) and (hState = 586)) or
								((vState = 96) and (hState = 587)) or
								((vState = 96) and (hState = 588)) or
								((vState = 96) and (hState = 593)) or
								((vState = 96) and (hState = 594)) or
								((vState = 96) and (hState = 596)) or
								((vState = 96) and (hState = 597)) or
								((vState = 96) and (hState = 598)) or
								((vState = 97) and (hState = 469)) or
								((vState = 97) and (hState = 470)) or
								((vState = 97) and (hState = 471)) or
								((vState = 97) and (hState = 472)) or
								((vState = 97) and (hState = 473)) or
								((vState = 97) and (hState = 474)) or
								((vState = 97) and (hState = 475)) or
								((vState = 97) and (hState = 476)) or
								((vState = 97) and (hState = 477)) or
								((vState = 97) and (hState = 478)) or
								((vState = 97) and (hState = 479)) or
								((vState = 97) and (hState = 480)) or
								((vState = 97) and (hState = 481)) or
								((vState = 97) and (hState = 482)) or
								((vState = 97) and (hState = 483)) or
								((vState = 97) and (hState = 484)) or
								((vState = 97) and (hState = 485)) or
								((vState = 97) and (hState = 486)) or
								((vState = 97) and (hState = 487)) or
								((vState = 97) and (hState = 488)) or
								((vState = 97) and (hState = 493)) or
								((vState = 97) and (hState = 494)) or
								((vState = 97) and (hState = 495)) or
								((vState = 97) and (hState = 499)) or
								((vState = 97) and (hState = 500)) or
								((vState = 97) and (hState = 501)) or
								((vState = 97) and (hState = 502)) or
								((vState = 97) and (hState = 503)) or
								((vState = 97) and (hState = 509)) or
								((vState = 97) and (hState = 510)) or
								((vState = 97) and (hState = 511)) or
								((vState = 97) and (hState = 517)) or
								((vState = 97) and (hState = 518)) or
								((vState = 97) and (hState = 519)) or
								((vState = 97) and (hState = 520)) or
								((vState = 97) and (hState = 521)) or
								((vState = 97) and (hState = 522)) or
								((vState = 97) and (hState = 526)) or
								((vState = 97) and (hState = 527)) or
								((vState = 97) and (hState = 528)) or
								((vState = 97) and (hState = 529)) or
								((vState = 97) and (hState = 535)) or
								((vState = 97) and (hState = 536)) or
								((vState = 97) and (hState = 539)) or
								((vState = 97) and (hState = 540)) or
								((vState = 97) and (hState = 541)) or
								((vState = 97) and (hState = 542)) or
								((vState = 97) and (hState = 543)) or
								((vState = 97) and (hState = 544)) or
								((vState = 97) and (hState = 546)) or
								((vState = 97) and (hState = 547)) or
								((vState = 97) and (hState = 548)) or
								((vState = 97) and (hState = 552)) or
								((vState = 97) and (hState = 553)) or
								((vState = 97) and (hState = 554)) or
								((vState = 97) and (hState = 555)) or
								((vState = 97) and (hState = 557)) or
								((vState = 97) and (hState = 558)) or
								((vState = 97) and (hState = 559)) or
								((vState = 97) and (hState = 560)) or
								((vState = 97) and (hState = 561)) or
								((vState = 97) and (hState = 562)) or
								((vState = 97) and (hState = 563)) or
								((vState = 97) and (hState = 564)) or
								((vState = 97) and (hState = 565)) or
								((vState = 97) and (hState = 566)) or
								((vState = 97) and (hState = 567)) or
								((vState = 97) and (hState = 568)) or
								((vState = 97) and (hState = 569)) or
								((vState = 97) and (hState = 571)) or
								((vState = 97) and (hState = 572)) or
								((vState = 97) and (hState = 573)) or
								((vState = 97) and (hState = 574)) or
								((vState = 97) and (hState = 575)) or
								((vState = 97) and (hState = 576)) or
								((vState = 97) and (hState = 577)) or
								((vState = 97) and (hState = 578)) or
								((vState = 97) and (hState = 581)) or
								((vState = 97) and (hState = 582)) or
								((vState = 97) and (hState = 583)) or
								((vState = 97) and (hState = 586)) or
								((vState = 97) and (hState = 587)) or
								((vState = 97) and (hState = 588)) or
								((vState = 97) and (hState = 592)) or
								((vState = 97) and (hState = 593)) or
								((vState = 97) and (hState = 594)) or
								((vState = 97) and (hState = 596)) or
								((vState = 97) and (hState = 597)) or
								((vState = 97) and (hState = 598)) or
								((vState = 98) and (hState = 468)) or
								((vState = 98) and (hState = 469)) or
								((vState = 98) and (hState = 470)) or
								((vState = 98) and (hState = 471)) or
								((vState = 98) and (hState = 472)) or
								((vState = 98) and (hState = 473)) or
								((vState = 98) and (hState = 474)) or
								((vState = 98) and (hState = 475)) or
								((vState = 98) and (hState = 476)) or
								((vState = 98) and (hState = 477)) or
								((vState = 98) and (hState = 478)) or
								((vState = 98) and (hState = 482)) or
								((vState = 98) and (hState = 483)) or
								((vState = 98) and (hState = 484)) or
								((vState = 98) and (hState = 485)) or
								((vState = 98) and (hState = 486)) or
								((vState = 98) and (hState = 487)) or
								((vState = 98) and (hState = 488)) or
								((vState = 98) and (hState = 489)) or
								((vState = 98) and (hState = 492)) or
								((vState = 98) and (hState = 494)) or
								((vState = 98) and (hState = 495)) or
								((vState = 98) and (hState = 499)) or
								((vState = 98) and (hState = 500)) or
								((vState = 98) and (hState = 501)) or
								((vState = 98) and (hState = 508)) or
								((vState = 98) and (hState = 509)) or
								((vState = 98) and (hState = 510)) or
								((vState = 98) and (hState = 517)) or
								((vState = 98) and (hState = 518)) or
								((vState = 98) and (hState = 519)) or
								((vState = 98) and (hState = 520)) or
								((vState = 98) and (hState = 521)) or
								((vState = 98) and (hState = 522)) or
								((vState = 98) and (hState = 523)) or
								((vState = 98) and (hState = 526)) or
								((vState = 98) and (hState = 527)) or
								((vState = 98) and (hState = 528)) or
								((vState = 98) and (hState = 529)) or
								((vState = 98) and (hState = 535)) or
								((vState = 98) and (hState = 536)) or
								((vState = 98) and (hState = 543)) or
								((vState = 98) and (hState = 544)) or
								((vState = 98) and (hState = 545)) or
								((vState = 98) and (hState = 546)) or
								((vState = 98) and (hState = 547)) or
								((vState = 98) and (hState = 548)) or
								((vState = 98) and (hState = 549)) or
								((vState = 98) and (hState = 551)) or
								((vState = 98) and (hState = 552)) or
								((vState = 98) and (hState = 553)) or
								((vState = 98) and (hState = 554)) or
								((vState = 98) and (hState = 555)) or
								((vState = 98) and (hState = 556)) or
								((vState = 98) and (hState = 557)) or
								((vState = 98) and (hState = 558)) or
								((vState = 98) and (hState = 559)) or
								((vState = 98) and (hState = 560)) or
								((vState = 98) and (hState = 561)) or
								((vState = 98) and (hState = 562)) or
								((vState = 98) and (hState = 563)) or
								((vState = 98) and (hState = 565)) or
								((vState = 98) and (hState = 566)) or
								((vState = 98) and (hState = 567)) or
								((vState = 98) and (hState = 568)) or
								((vState = 98) and (hState = 570)) or
								((vState = 98) and (hState = 571)) or
								((vState = 98) and (hState = 572)) or
								((vState = 98) and (hState = 573)) or
								((vState = 98) and (hState = 576)) or
								((vState = 98) and (hState = 577)) or
								((vState = 98) and (hState = 578)) or
								((vState = 98) and (hState = 580)) or
								((vState = 98) and (hState = 581)) or
								((vState = 98) and (hState = 582)) or
								((vState = 98) and (hState = 587)) or
								((vState = 98) and (hState = 588)) or
								((vState = 98) and (hState = 589)) or
								((vState = 98) and (hState = 592)) or
								((vState = 98) and (hState = 593)) or
								((vState = 98) and (hState = 596)) or
								((vState = 98) and (hState = 597)) or
								((vState = 98) and (hState = 598)) or
								((vState = 99) and (hState = 467)) or
								((vState = 99) and (hState = 468)) or
								((vState = 99) and (hState = 469)) or
								((vState = 99) and (hState = 470)) or
								((vState = 99) and (hState = 471)) or
								((vState = 99) and (hState = 472)) or
								((vState = 99) and (hState = 473)) or
								((vState = 99) and (hState = 474)) or
								((vState = 99) and (hState = 475)) or
								((vState = 99) and (hState = 482)) or
								((vState = 99) and (hState = 483)) or
								((vState = 99) and (hState = 484)) or
								((vState = 99) and (hState = 485)) or
								((vState = 99) and (hState = 486)) or
								((vState = 99) and (hState = 487)) or
								((vState = 99) and (hState = 488)) or
								((vState = 99) and (hState = 489)) or
								((vState = 99) and (hState = 492)) or
								((vState = 99) and (hState = 493)) or
								((vState = 99) and (hState = 495)) or
								((vState = 99) and (hState = 496)) or
								((vState = 99) and (hState = 498)) or
								((vState = 99) and (hState = 499)) or
								((vState = 99) and (hState = 500)) or
								((vState = 99) and (hState = 501)) or
								((vState = 99) and (hState = 507)) or
								((vState = 99) and (hState = 508)) or
								((vState = 99) and (hState = 509)) or
								((vState = 99) and (hState = 517)) or
								((vState = 99) and (hState = 518)) or
								((vState = 99) and (hState = 520)) or
								((vState = 99) and (hState = 521)) or
								((vState = 99) and (hState = 522)) or
								((vState = 99) and (hState = 523)) or
								((vState = 99) and (hState = 524)) or
								((vState = 99) and (hState = 525)) or
								((vState = 99) and (hState = 526)) or
								((vState = 99) and (hState = 535)) or
								((vState = 99) and (hState = 536)) or
								((vState = 99) and (hState = 544)) or
								((vState = 99) and (hState = 545)) or
								((vState = 99) and (hState = 546)) or
								((vState = 99) and (hState = 548)) or
								((vState = 99) and (hState = 549)) or
								((vState = 99) and (hState = 550)) or
								((vState = 99) and (hState = 551)) or
								((vState = 99) and (hState = 552)) or
								((vState = 99) and (hState = 553)) or
								((vState = 99) and (hState = 554)) or
								((vState = 99) and (hState = 555)) or
								((vState = 99) and (hState = 556)) or
								((vState = 99) and (hState = 557)) or
								((vState = 99) and (hState = 558)) or
								((vState = 99) and (hState = 559)) or
								((vState = 99) and (hState = 560)) or
								((vState = 99) and (hState = 562)) or
								((vState = 99) and (hState = 563)) or
								((vState = 99) and (hState = 564)) or
								((vState = 99) and (hState = 565)) or
								((vState = 99) and (hState = 566)) or
								((vState = 99) and (hState = 567)) or
								((vState = 99) and (hState = 568)) or
								((vState = 99) and (hState = 569)) or
								((vState = 99) and (hState = 570)) or
								((vState = 99) and (hState = 571)) or
								((vState = 99) and (hState = 572)) or
								((vState = 99) and (hState = 577)) or
								((vState = 99) and (hState = 578)) or
								((vState = 99) and (hState = 579)) or
								((vState = 99) and (hState = 580)) or
								((vState = 99) and (hState = 581)) or
								((vState = 99) and (hState = 587)) or
								((vState = 99) and (hState = 588)) or
								((vState = 99) and (hState = 589)) or
								((vState = 99) and (hState = 590)) or
								((vState = 99) and (hState = 591)) or
								((vState = 99) and (hState = 592)) or
								((vState = 99) and (hState = 593)) or
								((vState = 99) and (hState = 596)) or
								((vState = 99) and (hState = 597)) or
								((vState = 99) and (hState = 598)) or
								((vState = 100) and (hState = 466)) or
								((vState = 100) and (hState = 467)) or
								((vState = 100) and (hState = 468)) or
								((vState = 100) and (hState = 469)) or
								((vState = 100) and (hState = 475)) or
								((vState = 100) and (hState = 476)) or
								((vState = 100) and (hState = 482)) or
								((vState = 100) and (hState = 483)) or
								((vState = 100) and (hState = 484)) or
								((vState = 100) and (hState = 485)) or
								((vState = 100) and (hState = 486)) or
								((vState = 100) and (hState = 487)) or
								((vState = 100) and (hState = 488)) or
								((vState = 100) and (hState = 489)) or
								((vState = 100) and (hState = 490)) or
								((vState = 100) and (hState = 491)) or
								((vState = 100) and (hState = 492)) or
								((vState = 100) and (hState = 493)) or
								((vState = 100) and (hState = 494)) or
								((vState = 100) and (hState = 495)) or
								((vState = 100) and (hState = 496)) or
								((vState = 100) and (hState = 497)) or
								((vState = 100) and (hState = 498)) or
								((vState = 100) and (hState = 500)) or
								((vState = 100) and (hState = 501)) or
								((vState = 100) and (hState = 507)) or
								((vState = 100) and (hState = 508)) or
								((vState = 100) and (hState = 516)) or
								((vState = 100) and (hState = 517)) or
								((vState = 100) and (hState = 518)) or
								((vState = 100) and (hState = 520)) or
								((vState = 100) and (hState = 521)) or
								((vState = 100) and (hState = 522)) or
								((vState = 100) and (hState = 523)) or
								((vState = 100) and (hState = 524)) or
								((vState = 100) and (hState = 525)) or
								((vState = 100) and (hState = 526)) or
								((vState = 100) and (hState = 534)) or
								((vState = 100) and (hState = 535)) or
								((vState = 100) and (hState = 536)) or
								((vState = 100) and (hState = 545)) or
								((vState = 100) and (hState = 546)) or
								((vState = 100) and (hState = 547)) or
								((vState = 100) and (hState = 548)) or
								((vState = 100) and (hState = 549)) or
								((vState = 100) and (hState = 550)) or
								((vState = 100) and (hState = 551)) or
								((vState = 100) and (hState = 555)) or
								((vState = 100) and (hState = 556)) or
								((vState = 100) and (hState = 557)) or
								((vState = 100) and (hState = 559)) or
								((vState = 100) and (hState = 560)) or
								((vState = 100) and (hState = 561)) or
								((vState = 100) and (hState = 562)) or
								((vState = 100) and (hState = 563)) or
								((vState = 100) and (hState = 564)) or
								((vState = 100) and (hState = 565)) or
								((vState = 100) and (hState = 566)) or
								((vState = 100) and (hState = 567)) or
								((vState = 100) and (hState = 568)) or
								((vState = 100) and (hState = 569)) or
								((vState = 100) and (hState = 570)) or
								((vState = 100) and (hState = 571)) or
								((vState = 100) and (hState = 572)) or
								((vState = 100) and (hState = 576)) or
								((vState = 100) and (hState = 577)) or
								((vState = 100) and (hState = 578)) or
								((vState = 100) and (hState = 579)) or
								((vState = 100) and (hState = 580)) or
								((vState = 100) and (hState = 581)) or
								((vState = 100) and (hState = 587)) or
								((vState = 100) and (hState = 588)) or
								((vState = 100) and (hState = 589)) or
								((vState = 100) and (hState = 590)) or
								((vState = 100) and (hState = 591)) or
								((vState = 100) and (hState = 592)) or
								((vState = 100) and (hState = 597)) or
								((vState = 100) and (hState = 598)) or
								((vState = 101) and (hState = 475)) or
								((vState = 101) and (hState = 476)) or
								((vState = 101) and (hState = 482)) or
								((vState = 101) and (hState = 483)) or
								((vState = 101) and (hState = 484)) or
								((vState = 101) and (hState = 485)) or
								((vState = 101) and (hState = 486)) or
								((vState = 101) and (hState = 487)) or
								((vState = 101) and (hState = 488)) or
								((vState = 101) and (hState = 489)) or
								((vState = 101) and (hState = 490)) or
								((vState = 101) and (hState = 491)) or
								((vState = 101) and (hState = 492)) or
								((vState = 101) and (hState = 493)) or
								((vState = 101) and (hState = 494)) or
								((vState = 101) and (hState = 495)) or
								((vState = 101) and (hState = 496)) or
								((vState = 101) and (hState = 497)) or
								((vState = 101) and (hState = 500)) or
								((vState = 101) and (hState = 501)) or
								((vState = 101) and (hState = 507)) or
								((vState = 101) and (hState = 508)) or
								((vState = 101) and (hState = 516)) or
								((vState = 101) and (hState = 517)) or
								((vState = 101) and (hState = 518)) or
								((vState = 101) and (hState = 519)) or
								((vState = 101) and (hState = 520)) or
								((vState = 101) and (hState = 521)) or
								((vState = 101) and (hState = 522)) or
								((vState = 101) and (hState = 523)) or
								((vState = 101) and (hState = 524)) or
								((vState = 101) and (hState = 525)) or
								((vState = 101) and (hState = 526)) or
								((vState = 101) and (hState = 527)) or
								((vState = 101) and (hState = 534)) or
								((vState = 101) and (hState = 535)) or
								((vState = 101) and (hState = 536)) or
								((vState = 101) and (hState = 544)) or
								((vState = 101) and (hState = 545)) or
								((vState = 101) and (hState = 546)) or
								((vState = 101) and (hState = 547)) or
								((vState = 101) and (hState = 548)) or
								((vState = 101) and (hState = 549)) or
								((vState = 101) and (hState = 550)) or
								((vState = 101) and (hState = 551)) or
								((vState = 101) and (hState = 555)) or
								((vState = 101) and (hState = 556)) or
								((vState = 101) and (hState = 560)) or
								((vState = 101) and (hState = 561)) or
								((vState = 101) and (hState = 562)) or
								((vState = 101) and (hState = 563)) or
								((vState = 101) and (hState = 564)) or
								((vState = 101) and (hState = 565)) or
								((vState = 101) and (hState = 566)) or
								((vState = 101) and (hState = 567)) or
								((vState = 101) and (hState = 568)) or
								((vState = 101) and (hState = 569)) or
								((vState = 101) and (hState = 570)) or
								((vState = 101) and (hState = 571)) or
								((vState = 101) and (hState = 575)) or
								((vState = 101) and (hState = 576)) or
								((vState = 101) and (hState = 577)) or
								((vState = 101) and (hState = 578)) or
								((vState = 101) and (hState = 579)) or
								((vState = 101) and (hState = 580)) or
								((vState = 101) and (hState = 587)) or
								((vState = 101) and (hState = 588)) or
								((vState = 101) and (hState = 591)) or
								((vState = 101) and (hState = 592)) or
								((vState = 101) and (hState = 597)) or
								((vState = 101) and (hState = 598)) or
								((vState = 102) and (hState = 476)) or
								((vState = 102) and (hState = 477)) or
								((vState = 102) and (hState = 483)) or
								((vState = 102) and (hState = 484)) or
								((vState = 102) and (hState = 485)) or
								((vState = 102) and (hState = 486)) or
								((vState = 102) and (hState = 487)) or
								((vState = 102) and (hState = 488)) or
								((vState = 102) and (hState = 489)) or
								((vState = 102) and (hState = 490)) or
								((vState = 102) and (hState = 491)) or
								((vState = 102) and (hState = 492)) or
								((vState = 102) and (hState = 493)) or
								((vState = 102) and (hState = 494)) or
								((vState = 102) and (hState = 495)) or
								((vState = 102) and (hState = 496)) or
								((vState = 102) and (hState = 497)) or
								((vState = 102) and (hState = 500)) or
								((vState = 102) and (hState = 501)) or
								((vState = 102) and (hState = 507)) or
								((vState = 102) and (hState = 508)) or
								((vState = 102) and (hState = 515)) or
								((vState = 102) and (hState = 516)) or
								((vState = 102) and (hState = 517)) or
								((vState = 102) and (hState = 518)) or
								((vState = 102) and (hState = 519)) or
								((vState = 102) and (hState = 520)) or
								((vState = 102) and (hState = 521)) or
								((vState = 102) and (hState = 522)) or
								((vState = 102) and (hState = 523)) or
								((vState = 102) and (hState = 524)) or
								((vState = 102) and (hState = 526)) or
								((vState = 102) and (hState = 527)) or
								((vState = 102) and (hState = 528)) or
								((vState = 102) and (hState = 534)) or
								((vState = 102) and (hState = 535)) or
								((vState = 102) and (hState = 536)) or
								((vState = 102) and (hState = 537)) or
								((vState = 102) and (hState = 538)) or
								((vState = 102) and (hState = 539)) or
								((vState = 102) and (hState = 540)) or
								((vState = 102) and (hState = 544)) or
								((vState = 102) and (hState = 545)) or
								((vState = 102) and (hState = 548)) or
								((vState = 102) and (hState = 549)) or
								((vState = 102) and (hState = 550)) or
								((vState = 102) and (hState = 551)) or
								((vState = 102) and (hState = 552)) or
								((vState = 102) and (hState = 555)) or
								((vState = 102) and (hState = 556)) or
								((vState = 102) and (hState = 560)) or
								((vState = 102) and (hState = 561)) or
								((vState = 102) and (hState = 562)) or
								((vState = 102) and (hState = 563)) or
								((vState = 102) and (hState = 564)) or
								((vState = 102) and (hState = 565)) or
								((vState = 102) and (hState = 566)) or
								((vState = 102) and (hState = 567)) or
								((vState = 102) and (hState = 568)) or
								((vState = 102) and (hState = 569)) or
								((vState = 102) and (hState = 570)) or
								((vState = 102) and (hState = 571)) or
								((vState = 102) and (hState = 574)) or
								((vState = 102) and (hState = 575)) or
								((vState = 102) and (hState = 576)) or
								((vState = 102) and (hState = 577)) or
								((vState = 102) and (hState = 579)) or
								((vState = 102) and (hState = 580)) or
								((vState = 102) and (hState = 588)) or
								((vState = 102) and (hState = 591)) or
								((vState = 102) and (hState = 592)) or
								((vState = 102) and (hState = 593)) or
								((vState = 102) and (hState = 596)) or
								((vState = 102) and (hState = 597)) or
								((vState = 102) and (hState = 598)) or
								((vState = 103) and (hState = 476)) or
								((vState = 103) and (hState = 477)) or
								((vState = 103) and (hState = 478)) or
								((vState = 103) and (hState = 483)) or
								((vState = 103) and (hState = 484)) or
								((vState = 103) and (hState = 485)) or
								((vState = 103) and (hState = 486)) or
								((vState = 103) and (hState = 489)) or
								((vState = 103) and (hState = 490)) or
								((vState = 103) and (hState = 491)) or
								((vState = 103) and (hState = 492)) or
								((vState = 103) and (hState = 493)) or
								((vState = 103) and (hState = 494)) or
								((vState = 103) and (hState = 495)) or
								((vState = 103) and (hState = 496)) or
								((vState = 103) and (hState = 497)) or
								((vState = 103) and (hState = 498)) or
								((vState = 103) and (hState = 499)) or
								((vState = 103) and (hState = 500)) or
								((vState = 103) and (hState = 501)) or
								((vState = 103) and (hState = 507)) or
								((vState = 103) and (hState = 508)) or
								((vState = 103) and (hState = 514)) or
								((vState = 103) and (hState = 515)) or
								((vState = 103) and (hState = 516)) or
								((vState = 103) and (hState = 517)) or
								((vState = 103) and (hState = 518)) or
								((vState = 103) and (hState = 519)) or
								((vState = 103) and (hState = 520)) or
								((vState = 103) and (hState = 521)) or
								((vState = 103) and (hState = 522)) or
								((vState = 103) and (hState = 523)) or
								((vState = 103) and (hState = 524)) or
								((vState = 103) and (hState = 528)) or
								((vState = 103) and (hState = 529)) or
								((vState = 103) and (hState = 530)) or
								((vState = 103) and (hState = 531)) or
								((vState = 103) and (hState = 532)) or
								((vState = 103) and (hState = 533)) or
								((vState = 103) and (hState = 534)) or
								((vState = 103) and (hState = 535)) or
								((vState = 103) and (hState = 536)) or
								((vState = 103) and (hState = 537)) or
								((vState = 103) and (hState = 538)) or
								((vState = 103) and (hState = 539)) or
								((vState = 103) and (hState = 540)) or
								((vState = 103) and (hState = 541)) or
								((vState = 103) and (hState = 542)) or
								((vState = 103) and (hState = 543)) or
								((vState = 103) and (hState = 544)) or
								((vState = 103) and (hState = 545)) or
								((vState = 103) and (hState = 549)) or
								((vState = 103) and (hState = 550)) or
								((vState = 103) and (hState = 551)) or
								((vState = 103) and (hState = 552)) or
								((vState = 103) and (hState = 554)) or
								((vState = 103) and (hState = 555)) or
								((vState = 103) and (hState = 560)) or
								((vState = 103) and (hState = 561)) or
								((vState = 103) and (hState = 562)) or
								((vState = 103) and (hState = 563)) or
								((vState = 103) and (hState = 564)) or
								((vState = 103) and (hState = 565)) or
								((vState = 103) and (hState = 566)) or
								((vState = 103) and (hState = 567)) or
								((vState = 103) and (hState = 568)) or
								((vState = 103) and (hState = 569)) or
								((vState = 103) and (hState = 570)) or
								((vState = 103) and (hState = 571)) or
								((vState = 103) and (hState = 572)) or
								((vState = 103) and (hState = 573)) or
								((vState = 103) and (hState = 574)) or
								((vState = 103) and (hState = 575)) or
								((vState = 103) and (hState = 576)) or
								((vState = 103) and (hState = 577)) or
								((vState = 103) and (hState = 578)) or
								((vState = 103) and (hState = 579)) or
								((vState = 103) and (hState = 580)) or
								((vState = 103) and (hState = 581)) or
								((vState = 103) and (hState = 590)) or
								((vState = 103) and (hState = 591)) or
								((vState = 103) and (hState = 593)) or
								((vState = 103) and (hState = 594)) or
								((vState = 103) and (hState = 595)) or
								((vState = 103) and (hState = 596)) or
								((vState = 103) and (hState = 597)) or
								((vState = 103) and (hState = 598)) or
								((vState = 104) and (hState = 477)) or
								((vState = 104) and (hState = 478)) or
								((vState = 104) and (hState = 483)) or
								((vState = 104) and (hState = 484)) or
								((vState = 104) and (hState = 485)) or
								((vState = 104) and (hState = 486)) or
								((vState = 104) and (hState = 491)) or
								((vState = 104) and (hState = 492)) or
								((vState = 104) and (hState = 493)) or
								((vState = 104) and (hState = 494)) or
								((vState = 104) and (hState = 495)) or
								((vState = 104) and (hState = 496)) or
								((vState = 104) and (hState = 497)) or
								((vState = 104) and (hState = 498)) or
								((vState = 104) and (hState = 499)) or
								((vState = 104) and (hState = 500)) or
								((vState = 104) and (hState = 507)) or
								((vState = 104) and (hState = 508)) or
								((vState = 104) and (hState = 513)) or
								((vState = 104) and (hState = 514)) or
								((vState = 104) and (hState = 515)) or
								((vState = 104) and (hState = 517)) or
								((vState = 104) and (hState = 518)) or
								((vState = 104) and (hState = 519)) or
								((vState = 104) and (hState = 520)) or
								((vState = 104) and (hState = 521)) or
								((vState = 104) and (hState = 522)) or
								((vState = 104) and (hState = 523)) or
								((vState = 104) and (hState = 524)) or
								((vState = 104) and (hState = 529)) or
								((vState = 104) and (hState = 530)) or
								((vState = 104) and (hState = 531)) or
								((vState = 104) and (hState = 532)) or
								((vState = 104) and (hState = 533)) or
								((vState = 104) and (hState = 534)) or
								((vState = 104) and (hState = 535)) or
								((vState = 104) and (hState = 536)) or
								((vState = 104) and (hState = 537)) or
								((vState = 104) and (hState = 538)) or
								((vState = 104) and (hState = 539)) or
								((vState = 104) and (hState = 540)) or
								((vState = 104) and (hState = 541)) or
								((vState = 104) and (hState = 542)) or
								((vState = 104) and (hState = 543)) or
								((vState = 104) and (hState = 544)) or
								((vState = 104) and (hState = 545)) or
								((vState = 104) and (hState = 546)) or
								((vState = 104) and (hState = 547)) or
								((vState = 104) and (hState = 548)) or
								((vState = 104) and (hState = 550)) or
								((vState = 104) and (hState = 551)) or
								((vState = 104) and (hState = 552)) or
								((vState = 104) and (hState = 553)) or
								((vState = 104) and (hState = 554)) or
								((vState = 104) and (hState = 555)) or
								((vState = 104) and (hState = 560)) or
								((vState = 104) and (hState = 561)) or
								((vState = 104) and (hState = 562)) or
								((vState = 104) and (hState = 563)) or
								((vState = 104) and (hState = 564)) or
								((vState = 104) and (hState = 565)) or
								((vState = 104) and (hState = 566)) or
								((vState = 104) and (hState = 567)) or
								((vState = 104) and (hState = 568)) or
								((vState = 104) and (hState = 569)) or
								((vState = 104) and (hState = 570)) or
								((vState = 104) and (hState = 571)) or
								((vState = 104) and (hState = 572)) or
								((vState = 104) and (hState = 573)) or
								((vState = 104) and (hState = 574)) or
								((vState = 104) and (hState = 575)) or
								((vState = 104) and (hState = 576)) or
								((vState = 104) and (hState = 577)) or
								((vState = 104) and (hState = 578)) or
								((vState = 104) and (hState = 579)) or
								((vState = 104) and (hState = 580)) or
								((vState = 104) and (hState = 581)) or
								((vState = 104) and (hState = 582)) or
								((vState = 104) and (hState = 590)) or
								((vState = 104) and (hState = 591)) or
								((vState = 104) and (hState = 594)) or
								((vState = 104) and (hState = 595)) or
								((vState = 104) and (hState = 596)) or
								((vState = 104) and (hState = 597)) or
								((vState = 105) and (hState = 478)) or
								((vState = 105) and (hState = 479)) or
								((vState = 105) and (hState = 483)) or
								((vState = 105) and (hState = 484)) or
								((vState = 105) and (hState = 485)) or
								((vState = 105) and (hState = 486)) or
								((vState = 105) and (hState = 492)) or
								((vState = 105) and (hState = 493)) or
								((vState = 105) and (hState = 495)) or
								((vState = 105) and (hState = 496)) or
								((vState = 105) and (hState = 497)) or
								((vState = 105) and (hState = 498)) or
								((vState = 105) and (hState = 499)) or
								((vState = 105) and (hState = 500)) or
								((vState = 105) and (hState = 501)) or
								((vState = 105) and (hState = 507)) or
								((vState = 105) and (hState = 508)) or
								((vState = 105) and (hState = 513)) or
								((vState = 105) and (hState = 514)) or
								((vState = 105) and (hState = 517)) or
								((vState = 105) and (hState = 518)) or
								((vState = 105) and (hState = 519)) or
								((vState = 105) and (hState = 520)) or
								((vState = 105) and (hState = 521)) or
								((vState = 105) and (hState = 522)) or
								((vState = 105) and (hState = 524)) or
								((vState = 105) and (hState = 525)) or
								((vState = 105) and (hState = 531)) or
								((vState = 105) and (hState = 532)) or
								((vState = 105) and (hState = 533)) or
								((vState = 105) and (hState = 534)) or
								((vState = 105) and (hState = 542)) or
								((vState = 105) and (hState = 543)) or
								((vState = 105) and (hState = 544)) or
								((vState = 105) and (hState = 545)) or
								((vState = 105) and (hState = 546)) or
								((vState = 105) and (hState = 547)) or
								((vState = 105) and (hState = 548)) or
								((vState = 105) and (hState = 549)) or
								((vState = 105) and (hState = 550)) or
								((vState = 105) and (hState = 551)) or
								((vState = 105) and (hState = 552)) or
								((vState = 105) and (hState = 553)) or
								((vState = 105) and (hState = 554)) or
								((vState = 105) and (hState = 559)) or
								((vState = 105) and (hState = 560)) or
								((vState = 105) and (hState = 563)) or
								((vState = 105) and (hState = 564)) or
								((vState = 105) and (hState = 565)) or
								((vState = 105) and (hState = 569)) or
								((vState = 105) and (hState = 570)) or
								((vState = 105) and (hState = 571)) or
								((vState = 105) and (hState = 572)) or
								((vState = 105) and (hState = 573)) or
								((vState = 105) and (hState = 574)) or
								((vState = 105) and (hState = 575)) or
								((vState = 105) and (hState = 576)) or
								((vState = 105) and (hState = 577)) or
								((vState = 105) and (hState = 578)) or
								((vState = 105) and (hState = 579)) or
								((vState = 105) and (hState = 580)) or
								((vState = 105) and (hState = 589)) or
								((vState = 105) and (hState = 590)) or
								((vState = 105) and (hState = 594)) or
								((vState = 105) and (hState = 595)) or
								((vState = 105) and (hState = 596)) or
								((vState = 105) and (hState = 597)) or
								((vState = 106) and (hState = 479)) or
								((vState = 106) and (hState = 480)) or
								((vState = 106) and (hState = 483)) or
								((vState = 106) and (hState = 484)) or
								((vState = 106) and (hState = 485)) or
								((vState = 106) and (hState = 486)) or
								((vState = 106) and (hState = 492)) or
								((vState = 106) and (hState = 493)) or
								((vState = 106) and (hState = 496)) or
								((vState = 106) and (hState = 497)) or
								((vState = 106) and (hState = 498)) or
								((vState = 106) and (hState = 499)) or
								((vState = 106) and (hState = 500)) or
								((vState = 106) and (hState = 501)) or
								((vState = 106) and (hState = 502)) or
								((vState = 106) and (hState = 503)) or
								((vState = 106) and (hState = 508)) or
								((vState = 106) and (hState = 512)) or
								((vState = 106) and (hState = 513)) or
								((vState = 106) and (hState = 516)) or
								((vState = 106) and (hState = 517)) or
								((vState = 106) and (hState = 518)) or
								((vState = 106) and (hState = 519)) or
								((vState = 106) and (hState = 520)) or
								((vState = 106) and (hState = 521)) or
								((vState = 106) and (hState = 522)) or
								((vState = 106) and (hState = 523)) or
								((vState = 106) and (hState = 524)) or
								((vState = 106) and (hState = 525)) or
								((vState = 106) and (hState = 530)) or
								((vState = 106) and (hState = 531)) or
								((vState = 106) and (hState = 532)) or
								((vState = 106) and (hState = 533)) or
								((vState = 106) and (hState = 534)) or
								((vState = 106) and (hState = 540)) or
								((vState = 106) and (hState = 541)) or
								((vState = 106) and (hState = 542)) or
								((vState = 106) and (hState = 543)) or
								((vState = 106) and (hState = 544)) or
								((vState = 106) and (hState = 545)) or
								((vState = 106) and (hState = 546)) or
								((vState = 106) and (hState = 547)) or
								((vState = 106) and (hState = 548)) or
								((vState = 106) and (hState = 549)) or
								((vState = 106) and (hState = 550)) or
								((vState = 106) and (hState = 551)) or
								((vState = 106) and (hState = 552)) or
								((vState = 106) and (hState = 553)) or
								((vState = 106) and (hState = 554)) or
								((vState = 106) and (hState = 555)) or
								((vState = 106) and (hState = 558)) or
								((vState = 106) and (hState = 559)) or
								((vState = 106) and (hState = 560)) or
								((vState = 106) and (hState = 564)) or
								((vState = 106) and (hState = 565)) or
								((vState = 106) and (hState = 567)) or
								((vState = 106) and (hState = 568)) or
								((vState = 106) and (hState = 569)) or
								((vState = 106) and (hState = 570)) or
								((vState = 106) and (hState = 571)) or
								((vState = 106) and (hState = 572)) or
								((vState = 106) and (hState = 573)) or
								((vState = 106) and (hState = 574)) or
								((vState = 106) and (hState = 575)) or
								((vState = 106) and (hState = 576)) or
								((vState = 106) and (hState = 577)) or
								((vState = 106) and (hState = 578)) or
								((vState = 106) and (hState = 588)) or
								((vState = 106) and (hState = 589)) or
								((vState = 106) and (hState = 590)) or
								((vState = 106) and (hState = 594)) or
								((vState = 106) and (hState = 595)) or
								((vState = 106) and (hState = 596)) or
								((vState = 106) and (hState = 597)) or
								((vState = 107) and (hState = 479)) or
								((vState = 107) and (hState = 480)) or
								((vState = 107) and (hState = 481)) or
								((vState = 107) and (hState = 484)) or
								((vState = 107) and (hState = 485)) or
								((vState = 107) and (hState = 492)) or
								((vState = 107) and (hState = 493)) or
								((vState = 107) and (hState = 497)) or
								((vState = 107) and (hState = 498)) or
								((vState = 107) and (hState = 499)) or
								((vState = 107) and (hState = 500)) or
								((vState = 107) and (hState = 501)) or
								((vState = 107) and (hState = 502)) or
								((vState = 107) and (hState = 503)) or
								((vState = 107) and (hState = 504)) or
								((vState = 107) and (hState = 505)) or
								((vState = 107) and (hState = 508)) or
								((vState = 107) and (hState = 509)) or
								((vState = 107) and (hState = 512)) or
								((vState = 107) and (hState = 513)) or
								((vState = 107) and (hState = 516)) or
								((vState = 107) and (hState = 517)) or
								((vState = 107) and (hState = 518)) or
								((vState = 107) and (hState = 519)) or
								((vState = 107) and (hState = 520)) or
								((vState = 107) and (hState = 521)) or
								((vState = 107) and (hState = 522)) or
								((vState = 107) and (hState = 523)) or
								((vState = 107) and (hState = 524)) or
								((vState = 107) and (hState = 525)) or
								((vState = 107) and (hState = 529)) or
								((vState = 107) and (hState = 530)) or
								((vState = 107) and (hState = 533)) or
								((vState = 107) and (hState = 534)) or
								((vState = 107) and (hState = 537)) or
								((vState = 107) and (hState = 538)) or
								((vState = 107) and (hState = 539)) or
								((vState = 107) and (hState = 540)) or
								((vState = 107) and (hState = 541)) or
								((vState = 107) and (hState = 542)) or
								((vState = 107) and (hState = 543)) or
								((vState = 107) and (hState = 544)) or
								((vState = 107) and (hState = 545)) or
								((vState = 107) and (hState = 546)) or
								((vState = 107) and (hState = 547)) or
								((vState = 107) and (hState = 548)) or
								((vState = 107) and (hState = 549)) or
								((vState = 107) and (hState = 550)) or
								((vState = 107) and (hState = 551)) or
								((vState = 107) and (hState = 552)) or
								((vState = 107) and (hState = 553)) or
								((vState = 107) and (hState = 554)) or
								((vState = 107) and (hState = 555)) or
								((vState = 107) and (hState = 556)) or
								((vState = 107) and (hState = 557)) or
								((vState = 107) and (hState = 558)) or
								((vState = 107) and (hState = 559)) or
								((vState = 107) and (hState = 564)) or
								((vState = 107) and (hState = 565)) or
								((vState = 107) and (hState = 566)) or
								((vState = 107) and (hState = 567)) or
								((vState = 107) and (hState = 568)) or
								((vState = 107) and (hState = 569)) or
								((vState = 107) and (hState = 570)) or
								((vState = 107) and (hState = 571)) or
								((vState = 107) and (hState = 572)) or
								((vState = 107) and (hState = 573)) or
								((vState = 107) and (hState = 574)) or
								((vState = 107) and (hState = 577)) or
								((vState = 107) and (hState = 578)) or
								((vState = 107) and (hState = 588)) or
								((vState = 107) and (hState = 589)) or
								((vState = 107) and (hState = 593)) or
								((vState = 107) and (hState = 594)) or
								((vState = 107) and (hState = 595)) or
								((vState = 107) and (hState = 596)) or
								((vState = 107) and (hState = 597)) or
								((vState = 107) and (hState = 598)) or
								((vState = 108) and (hState = 480)) or
								((vState = 108) and (hState = 481)) or
								((vState = 108) and (hState = 484)) or
								((vState = 108) and (hState = 485)) or
								((vState = 108) and (hState = 492)) or
								((vState = 108) and (hState = 493)) or
								((vState = 108) and (hState = 498)) or
								((vState = 108) and (hState = 499)) or
								((vState = 108) and (hState = 500)) or
								((vState = 108) and (hState = 501)) or
								((vState = 108) and (hState = 504)) or
								((vState = 108) and (hState = 505)) or
								((vState = 108) and (hState = 506)) or
								((vState = 108) and (hState = 507)) or
								((vState = 108) and (hState = 508)) or
								((vState = 108) and (hState = 509)) or
								((vState = 108) and (hState = 511)) or
								((vState = 108) and (hState = 512)) or
								((vState = 108) and (hState = 516)) or
								((vState = 108) and (hState = 517)) or
								((vState = 108) and (hState = 518)) or
								((vState = 108) and (hState = 519)) or
								((vState = 108) and (hState = 520)) or
								((vState = 108) and (hState = 523)) or
								((vState = 108) and (hState = 524)) or
								((vState = 108) and (hState = 525)) or
								((vState = 108) and (hState = 526)) or
								((vState = 108) and (hState = 528)) or
								((vState = 108) and (hState = 529)) or
								((vState = 108) and (hState = 533)) or
								((vState = 108) and (hState = 534)) or
								((vState = 108) and (hState = 536)) or
								((vState = 108) and (hState = 537)) or
								((vState = 108) and (hState = 540)) or
								((vState = 108) and (hState = 541)) or
								((vState = 108) and (hState = 542)) or
								((vState = 108) and (hState = 544)) or
								((vState = 108) and (hState = 545)) or
								((vState = 108) and (hState = 546)) or
								((vState = 108) and (hState = 552)) or
								((vState = 108) and (hState = 553)) or
								((vState = 108) and (hState = 554)) or
								((vState = 108) and (hState = 555)) or
								((vState = 108) and (hState = 556)) or
								((vState = 108) and (hState = 557)) or
								((vState = 108) and (hState = 558)) or
								((vState = 108) and (hState = 559)) or
								((vState = 108) and (hState = 560)) or
								((vState = 108) and (hState = 561)) or
								((vState = 108) and (hState = 562)) or
								((vState = 108) and (hState = 563)) or
								((vState = 108) and (hState = 564)) or
								((vState = 108) and (hState = 565)) or
								((vState = 108) and (hState = 566)) or
								((vState = 108) and (hState = 567)) or
								((vState = 108) and (hState = 568)) or
								((vState = 108) and (hState = 569)) or
								((vState = 108) and (hState = 570)) or
								((vState = 108) and (hState = 571)) or
								((vState = 108) and (hState = 572)) or
								((vState = 108) and (hState = 573)) or
								((vState = 108) and (hState = 574)) or
								((vState = 108) and (hState = 575)) or
								((vState = 108) and (hState = 576)) or
								((vState = 108) and (hState = 577)) or
								((vState = 108) and (hState = 587)) or
								((vState = 108) and (hState = 588)) or
								((vState = 108) and (hState = 592)) or
								((vState = 108) and (hState = 593)) or
								((vState = 108) and (hState = 595)) or
								((vState = 108) and (hState = 596)) or
								((vState = 108) and (hState = 598)) or
								((vState = 108) and (hState = 599)) or
								((vState = 109) and (hState = 481)) or
								((vState = 109) and (hState = 482)) or
								((vState = 109) and (hState = 484)) or
								((vState = 109) and (hState = 485)) or
								((vState = 109) and (hState = 492)) or
								((vState = 109) and (hState = 493)) or
								((vState = 109) and (hState = 498)) or
								((vState = 109) and (hState = 499)) or
								((vState = 109) and (hState = 500)) or
								((vState = 109) and (hState = 501)) or
								((vState = 109) and (hState = 506)) or
								((vState = 109) and (hState = 507)) or
								((vState = 109) and (hState = 508)) or
								((vState = 109) and (hState = 509)) or
								((vState = 109) and (hState = 510)) or
								((vState = 109) and (hState = 511)) or
								((vState = 109) and (hState = 512)) or
								((vState = 109) and (hState = 516)) or
								((vState = 109) and (hState = 517)) or
								((vState = 109) and (hState = 518)) or
								((vState = 109) and (hState = 519)) or
								((vState = 109) and (hState = 524)) or
								((vState = 109) and (hState = 525)) or
								((vState = 109) and (hState = 526)) or
								((vState = 109) and (hState = 527)) or
								((vState = 109) and (hState = 528)) or
								((vState = 109) and (hState = 533)) or
								((vState = 109) and (hState = 534)) or
								((vState = 109) and (hState = 535)) or
								((vState = 109) and (hState = 536)) or
								((vState = 109) and (hState = 540)) or
								((vState = 109) and (hState = 541)) or
								((vState = 109) and (hState = 542)) or
								((vState = 109) and (hState = 543)) or
								((vState = 109) and (hState = 544)) or
								((vState = 109) and (hState = 545)) or
								((vState = 109) and (hState = 546)) or
								((vState = 109) and (hState = 547)) or
								((vState = 109) and (hState = 551)) or
								((vState = 109) and (hState = 552)) or
								((vState = 109) and (hState = 555)) or
								((vState = 109) and (hState = 556)) or
								((vState = 109) and (hState = 557)) or
								((vState = 109) and (hState = 558)) or
								((vState = 109) and (hState = 561)) or
								((vState = 109) and (hState = 562)) or
								((vState = 109) and (hState = 563)) or
								((vState = 109) and (hState = 564)) or
								((vState = 109) and (hState = 565)) or
								((vState = 109) and (hState = 566)) or
								((vState = 109) and (hState = 567)) or
								((vState = 109) and (hState = 568)) or
								((vState = 109) and (hState = 569)) or
								((vState = 109) and (hState = 570)) or
								((vState = 109) and (hState = 571)) or
								((vState = 109) and (hState = 572)) or
								((vState = 109) and (hState = 573)) or
								((vState = 109) and (hState = 574)) or
								((vState = 109) and (hState = 575)) or
								((vState = 109) and (hState = 576)) or
								((vState = 109) and (hState = 577)) or
								((vState = 109) and (hState = 587)) or
								((vState = 109) and (hState = 588)) or
								((vState = 109) and (hState = 591)) or
								((vState = 109) and (hState = 592)) or
								((vState = 109) and (hState = 593)) or
								((vState = 109) and (hState = 595)) or
								((vState = 109) and (hState = 596)) or
								((vState = 109) and (hState = 599)) or
								((vState = 110) and (hState = 482)) or
								((vState = 110) and (hState = 483)) or
								((vState = 110) and (hState = 484)) or
								((vState = 110) and (hState = 485)) or
								((vState = 110) and (hState = 492)) or
								((vState = 110) and (hState = 493)) or
								((vState = 110) and (hState = 497)) or
								((vState = 110) and (hState = 498)) or
								((vState = 110) and (hState = 499)) or
								((vState = 110) and (hState = 500)) or
								((vState = 110) and (hState = 501)) or
								((vState = 110) and (hState = 502)) or
								((vState = 110) and (hState = 508)) or
								((vState = 110) and (hState = 509)) or
								((vState = 110) and (hState = 510)) or
								((vState = 110) and (hState = 511)) or
								((vState = 110) and (hState = 512)) or
								((vState = 110) and (hState = 516)) or
								((vState = 110) and (hState = 517)) or
								((vState = 110) and (hState = 518)) or
								((vState = 110) and (hState = 525)) or
								((vState = 110) and (hState = 526)) or
								((vState = 110) and (hState = 527)) or
								((vState = 110) and (hState = 528)) or
								((vState = 110) and (hState = 532)) or
								((vState = 110) and (hState = 533)) or
								((vState = 110) and (hState = 534)) or
								((vState = 110) and (hState = 535)) or
								((vState = 110) and (hState = 540)) or
								((vState = 110) and (hState = 541)) or
								((vState = 110) and (hState = 542)) or
								((vState = 110) and (hState = 543)) or
								((vState = 110) and (hState = 544)) or
								((vState = 110) and (hState = 545)) or
								((vState = 110) and (hState = 546)) or
								((vState = 110) and (hState = 547)) or
								((vState = 110) and (hState = 548)) or
								((vState = 110) and (hState = 549)) or
								((vState = 110) and (hState = 550)) or
								((vState = 110) and (hState = 551)) or
								((vState = 110) and (hState = 552)) or
								((vState = 110) and (hState = 554)) or
								((vState = 110) and (hState = 555)) or
								((vState = 110) and (hState = 556)) or
								((vState = 110) and (hState = 557)) or
								((vState = 110) and (hState = 558)) or
								((vState = 110) and (hState = 565)) or
								((vState = 110) and (hState = 566)) or
								((vState = 110) and (hState = 567)) or
								((vState = 110) and (hState = 568)) or
								((vState = 110) and (hState = 569)) or
								((vState = 110) and (hState = 570)) or
								((vState = 110) and (hState = 574)) or
								((vState = 110) and (hState = 575)) or
								((vState = 110) and (hState = 576)) or
								((vState = 110) and (hState = 586)) or
								((vState = 110) and (hState = 587)) or
								((vState = 110) and (hState = 590)) or
								((vState = 110) and (hState = 591)) or
								((vState = 110) and (hState = 592)) or
								((vState = 110) and (hState = 595)) or
								((vState = 110) and (hState = 596)) or
								((vState = 111) and (hState = 483)) or
								((vState = 111) and (hState = 484)) or
								((vState = 111) and (hState = 485)) or
								((vState = 111) and (hState = 492)) or
								((vState = 111) and (hState = 493)) or
								((vState = 111) and (hState = 497)) or
								((vState = 111) and (hState = 498)) or
								((vState = 111) and (hState = 500)) or
								((vState = 111) and (hState = 501)) or
								((vState = 111) and (hState = 502)) or
								((vState = 111) and (hState = 508)) or
								((vState = 111) and (hState = 509)) or
								((vState = 111) and (hState = 510)) or
								((vState = 111) and (hState = 511)) or
								((vState = 111) and (hState = 512)) or
								((vState = 111) and (hState = 513)) or
								((vState = 111) and (hState = 514)) or
								((vState = 111) and (hState = 515)) or
								((vState = 111) and (hState = 516)) or
								((vState = 111) and (hState = 517)) or
								((vState = 111) and (hState = 518)) or
								((vState = 111) and (hState = 524)) or
								((vState = 111) and (hState = 525)) or
								((vState = 111) and (hState = 526)) or
								((vState = 111) and (hState = 527)) or
								((vState = 111) and (hState = 528)) or
								((vState = 111) and (hState = 532)) or
								((vState = 111) and (hState = 533)) or
								((vState = 111) and (hState = 534)) or
								((vState = 111) and (hState = 539)) or
								((vState = 111) and (hState = 540)) or
								((vState = 111) and (hState = 541)) or
								((vState = 111) and (hState = 542)) or
								((vState = 111) and (hState = 543)) or
								((vState = 111) and (hState = 544)) or
								((vState = 111) and (hState = 545)) or
								((vState = 111) and (hState = 546)) or
								((vState = 111) and (hState = 549)) or
								((vState = 111) and (hState = 550)) or
								((vState = 111) and (hState = 551)) or
								((vState = 111) and (hState = 552)) or
								((vState = 111) and (hState = 553)) or
								((vState = 111) and (hState = 554)) or
								((vState = 111) and (hState = 558)) or
								((vState = 111) and (hState = 559)) or
								((vState = 111) and (hState = 565)) or
								((vState = 111) and (hState = 566)) or
								((vState = 111) and (hState = 567)) or
								((vState = 111) and (hState = 568)) or
								((vState = 111) and (hState = 569)) or
								((vState = 111) and (hState = 575)) or
								((vState = 111) and (hState = 576)) or
								((vState = 111) and (hState = 585)) or
								((vState = 111) and (hState = 586)) or
								((vState = 111) and (hState = 589)) or
								((vState = 111) and (hState = 590)) or
								((vState = 111) and (hState = 591)) or
								((vState = 111) and (hState = 595)) or
								((vState = 111) and (hState = 596)) or
								((vState = 112) and (hState = 483)) or
								((vState = 112) and (hState = 484)) or
								((vState = 112) and (hState = 485)) or
								((vState = 112) and (hState = 492)) or
								((vState = 112) and (hState = 493)) or
								((vState = 112) and (hState = 494)) or
								((vState = 112) and (hState = 495)) or
								((vState = 112) and (hState = 496)) or
								((vState = 112) and (hState = 497)) or
								((vState = 112) and (hState = 498)) or
								((vState = 112) and (hState = 499)) or
								((vState = 112) and (hState = 500)) or
								((vState = 112) and (hState = 501)) or
								((vState = 112) and (hState = 502)) or
								((vState = 112) and (hState = 503)) or
								((vState = 112) and (hState = 508)) or
								((vState = 112) and (hState = 509)) or
								((vState = 112) and (hState = 510)) or
								((vState = 112) and (hState = 513)) or
								((vState = 112) and (hState = 514)) or
								((vState = 112) and (hState = 515)) or
								((vState = 112) and (hState = 516)) or
								((vState = 112) and (hState = 517)) or
								((vState = 112) and (hState = 524)) or
								((vState = 112) and (hState = 525)) or
								((vState = 112) and (hState = 526)) or
								((vState = 112) and (hState = 527)) or
								((vState = 112) and (hState = 528)) or
								((vState = 112) and (hState = 529)) or
								((vState = 112) and (hState = 530)) or
								((vState = 112) and (hState = 532)) or
								((vState = 112) and (hState = 533)) or
								((vState = 112) and (hState = 534)) or
								((vState = 112) and (hState = 535)) or
								((vState = 112) and (hState = 536)) or
								((vState = 112) and (hState = 537)) or
								((vState = 112) and (hState = 538)) or
								((vState = 112) and (hState = 539)) or
								((vState = 112) and (hState = 540)) or
								((vState = 112) and (hState = 541)) or
								((vState = 112) and (hState = 545)) or
								((vState = 112) and (hState = 546)) or
								((vState = 112) and (hState = 547)) or
								((vState = 112) and (hState = 550)) or
								((vState = 112) and (hState = 551)) or
								((vState = 112) and (hState = 552)) or
								((vState = 112) and (hState = 553)) or
								((vState = 112) and (hState = 554)) or
								((vState = 112) and (hState = 555)) or
								((vState = 112) and (hState = 556)) or
								((vState = 112) and (hState = 557)) or
								((vState = 112) and (hState = 558)) or
								((vState = 112) and (hState = 559)) or
								((vState = 112) and (hState = 560)) or
								((vState = 112) and (hState = 565)) or
								((vState = 112) and (hState = 566)) or
								((vState = 112) and (hState = 567)) or
								((vState = 112) and (hState = 568)) or
								((vState = 112) and (hState = 569)) or
								((vState = 112) and (hState = 576)) or
								((vState = 112) and (hState = 577)) or
								((vState = 112) and (hState = 583)) or
								((vState = 112) and (hState = 584)) or
								((vState = 112) and (hState = 585)) or
								((vState = 112) and (hState = 586)) or
								((vState = 112) and (hState = 588)) or
								((vState = 112) and (hState = 589)) or
								((vState = 112) and (hState = 590)) or
								((vState = 112) and (hState = 595)) or
								((vState = 112) and (hState = 596)) or
								((vState = 113) and (hState = 484)) or
								((vState = 113) and (hState = 485)) or
								((vState = 113) and (hState = 495)) or
								((vState = 113) and (hState = 496)) or
								((vState = 113) and (hState = 497)) or
								((vState = 113) and (hState = 498)) or
								((vState = 113) and (hState = 499)) or
								((vState = 113) and (hState = 500)) or
								((vState = 113) and (hState = 501)) or
								((vState = 113) and (hState = 502)) or
								((vState = 113) and (hState = 503)) or
								((vState = 113) and (hState = 509)) or
								((vState = 113) and (hState = 514)) or
								((vState = 113) and (hState = 515)) or
								((vState = 113) and (hState = 516)) or
								((vState = 113) and (hState = 517)) or
								((vState = 113) and (hState = 518)) or
								((vState = 113) and (hState = 522)) or
								((vState = 113) and (hState = 523)) or
								((vState = 113) and (hState = 524)) or
								((vState = 113) and (hState = 525)) or
								((vState = 113) and (hState = 526)) or
								((vState = 113) and (hState = 527)) or
								((vState = 113) and (hState = 529)) or
								((vState = 113) and (hState = 530)) or
								((vState = 113) and (hState = 531)) or
								((vState = 113) and (hState = 532)) or
								((vState = 113) and (hState = 533)) or
								((vState = 113) and (hState = 534)) or
								((vState = 113) and (hState = 535)) or
								((vState = 113) and (hState = 536)) or
								((vState = 113) and (hState = 537)) or
								((vState = 113) and (hState = 538)) or
								((vState = 113) and (hState = 539)) or
								((vState = 113) and (hState = 540)) or
								((vState = 113) and (hState = 546)) or
								((vState = 113) and (hState = 547)) or
								((vState = 113) and (hState = 548)) or
								((vState = 113) and (hState = 549)) or
								((vState = 113) and (hState = 550)) or
								((vState = 113) and (hState = 551)) or
								((vState = 113) and (hState = 552)) or
								((vState = 113) and (hState = 553)) or
								((vState = 113) and (hState = 554)) or
								((vState = 113) and (hState = 555)) or
								((vState = 113) and (hState = 556)) or
								((vState = 113) and (hState = 557)) or
								((vState = 113) and (hState = 558)) or
								((vState = 113) and (hState = 559)) or
								((vState = 113) and (hState = 560)) or
								((vState = 113) and (hState = 561)) or
								((vState = 113) and (hState = 564)) or
								((vState = 113) and (hState = 565)) or
								((vState = 113) and (hState = 566)) or
								((vState = 113) and (hState = 567)) or
								((vState = 113) and (hState = 568)) or
								((vState = 113) and (hState = 569)) or
								((vState = 113) and (hState = 570)) or
								((vState = 113) and (hState = 576)) or
								((vState = 113) and (hState = 577)) or
								((vState = 113) and (hState = 582)) or
								((vState = 113) and (hState = 583)) or
								((vState = 113) and (hState = 584)) or
								((vState = 113) and (hState = 585)) or
								((vState = 113) and (hState = 586)) or
								((vState = 113) and (hState = 588)) or
								((vState = 113) and (hState = 589)) or
								((vState = 113) and (hState = 594)) or
								((vState = 113) and (hState = 595)) or
								((vState = 114) and (hState = 485)) or
								((vState = 114) and (hState = 486)) or
								((vState = 114) and (hState = 498)) or
								((vState = 114) and (hState = 499)) or
								((vState = 114) and (hState = 500)) or
								((vState = 114) and (hState = 501)) or
								((vState = 114) and (hState = 502)) or
								((vState = 114) and (hState = 503)) or
								((vState = 114) and (hState = 504)) or
								((vState = 114) and (hState = 514)) or
								((vState = 114) and (hState = 515)) or
								((vState = 114) and (hState = 516)) or
								((vState = 114) and (hState = 517)) or
								((vState = 114) and (hState = 518)) or
								((vState = 114) and (hState = 519)) or
								((vState = 114) and (hState = 520)) or
								((vState = 114) and (hState = 521)) or
								((vState = 114) and (hState = 522)) or
								((vState = 114) and (hState = 523)) or
								((vState = 114) and (hState = 526)) or
								((vState = 114) and (hState = 527)) or
								((vState = 114) and (hState = 530)) or
								((vState = 114) and (hState = 531)) or
								((vState = 114) and (hState = 532)) or
								((vState = 114) and (hState = 536)) or
								((vState = 114) and (hState = 537)) or
								((vState = 114) and (hState = 538)) or
								((vState = 114) and (hState = 539)) or
								((vState = 114) and (hState = 547)) or
								((vState = 114) and (hState = 548)) or
								((vState = 114) and (hState = 549)) or
								((vState = 114) and (hState = 550)) or
								((vState = 114) and (hState = 551)) or
								((vState = 114) and (hState = 558)) or
								((vState = 114) and (hState = 559)) or
								((vState = 114) and (hState = 560)) or
								((vState = 114) and (hState = 561)) or
								((vState = 114) and (hState = 562)) or
								((vState = 114) and (hState = 563)) or
								((vState = 114) and (hState = 564)) or
								((vState = 114) and (hState = 565)) or
								((vState = 114) and (hState = 566)) or
								((vState = 114) and (hState = 567)) or
								((vState = 114) and (hState = 568)) or
								((vState = 114) and (hState = 570)) or
								((vState = 114) and (hState = 571)) or
								((vState = 114) and (hState = 577)) or
								((vState = 114) and (hState = 580)) or
								((vState = 114) and (hState = 581)) or
								((vState = 114) and (hState = 582)) or
								((vState = 114) and (hState = 583)) or
								((vState = 114) and (hState = 584)) or
								((vState = 114) and (hState = 585)) or
								((vState = 114) and (hState = 586)) or
								((vState = 114) and (hState = 587)) or
								((vState = 114) and (hState = 588)) or
								((vState = 114) and (hState = 593)) or
								((vState = 114) and (hState = 594)) or
								((vState = 114) and (hState = 595)) or
								((vState = 115) and (hState = 486)) or
								((vState = 115) and (hState = 487)) or
								((vState = 115) and (hState = 500)) or
								((vState = 115) and (hState = 501)) or
								((vState = 115) and (hState = 502)) or
								((vState = 115) and (hState = 503)) or
								((vState = 115) and (hState = 504)) or
								((vState = 115) and (hState = 505)) or
								((vState = 115) and (hState = 506)) or
								((vState = 115) and (hState = 507)) or
								((vState = 115) and (hState = 513)) or
								((vState = 115) and (hState = 514)) or
								((vState = 115) and (hState = 515)) or
								((vState = 115) and (hState = 516)) or
								((vState = 115) and (hState = 517)) or
								((vState = 115) and (hState = 519)) or
								((vState = 115) and (hState = 520)) or
								((vState = 115) and (hState = 521)) or
								((vState = 115) and (hState = 522)) or
								((vState = 115) and (hState = 526)) or
								((vState = 115) and (hState = 527)) or
								((vState = 115) and (hState = 529)) or
								((vState = 115) and (hState = 530)) or
								((vState = 115) and (hState = 531)) or
								((vState = 115) and (hState = 532)) or
								((vState = 115) and (hState = 533)) or
								((vState = 115) and (hState = 536)) or
								((vState = 115) and (hState = 537)) or
								((vState = 115) and (hState = 538)) or
								((vState = 115) and (hState = 548)) or
								((vState = 115) and (hState = 549)) or
								((vState = 115) and (hState = 550)) or
								((vState = 115) and (hState = 561)) or
								((vState = 115) and (hState = 562)) or
								((vState = 115) and (hState = 563)) or
								((vState = 115) and (hState = 566)) or
								((vState = 115) and (hState = 567)) or
								((vState = 115) and (hState = 570)) or
								((vState = 115) and (hState = 571)) or
								((vState = 115) and (hState = 572)) or
								((vState = 115) and (hState = 576)) or
								((vState = 115) and (hState = 577)) or
								((vState = 115) and (hState = 578)) or
								((vState = 115) and (hState = 579)) or
								((vState = 115) and (hState = 580)) or
								((vState = 115) and (hState = 581)) or
								((vState = 115) and (hState = 582)) or
								((vState = 115) and (hState = 583)) or
								((vState = 115) and (hState = 584)) or
								((vState = 115) and (hState = 585)) or
								((vState = 115) and (hState = 586)) or
								((vState = 115) and (hState = 587)) or
								((vState = 115) and (hState = 592)) or
								((vState = 115) and (hState = 593)) or
								((vState = 115) and (hState = 594)) or
								((vState = 115) and (hState = 595)) or
								((vState = 116) and (hState = 486)) or
								((vState = 116) and (hState = 487)) or
								((vState = 116) and (hState = 488)) or
								((vState = 116) and (hState = 490)) or
								((vState = 116) and (hState = 491)) or
								((vState = 116) and (hState = 492)) or
								((vState = 116) and (hState = 493)) or
								((vState = 116) and (hState = 494)) or
								((vState = 116) and (hState = 495)) or
								((vState = 116) and (hState = 496)) or
								((vState = 116) and (hState = 497)) or
								((vState = 116) and (hState = 498)) or
								((vState = 116) and (hState = 499)) or
								((vState = 116) and (hState = 500)) or
								((vState = 116) and (hState = 501)) or
								((vState = 116) and (hState = 502)) or
								((vState = 116) and (hState = 503)) or
								((vState = 116) and (hState = 504)) or
								((vState = 116) and (hState = 505)) or
								((vState = 116) and (hState = 506)) or
								((vState = 116) and (hState = 507)) or
								((vState = 116) and (hState = 508)) or
								((vState = 116) and (hState = 509)) or
								((vState = 116) and (hState = 512)) or
								((vState = 116) and (hState = 513)) or
								((vState = 116) and (hState = 514)) or
								((vState = 116) and (hState = 515)) or
								((vState = 116) and (hState = 516)) or
								((vState = 116) and (hState = 517)) or
								((vState = 116) and (hState = 524)) or
								((vState = 116) and (hState = 525)) or
								((vState = 116) and (hState = 526)) or
								((vState = 116) and (hState = 527)) or
								((vState = 116) and (hState = 528)) or
								((vState = 116) and (hState = 529)) or
								((vState = 116) and (hState = 533)) or
								((vState = 116) and (hState = 534)) or
								((vState = 116) and (hState = 535)) or
								((vState = 116) and (hState = 536)) or
								((vState = 116) and (hState = 537)) or
								((vState = 116) and (hState = 548)) or
								((vState = 116) and (hState = 549)) or
								((vState = 116) and (hState = 550)) or
								((vState = 116) and (hState = 560)) or
								((vState = 116) and (hState = 561)) or
								((vState = 116) and (hState = 562)) or
								((vState = 116) and (hState = 567)) or
								((vState = 116) and (hState = 569)) or
								((vState = 116) and (hState = 570)) or
								((vState = 116) and (hState = 571)) or
								((vState = 116) and (hState = 576)) or
								((vState = 116) and (hState = 577)) or
								((vState = 116) and (hState = 578)) or
								((vState = 116) and (hState = 579)) or
								((vState = 116) and (hState = 580)) or
								((vState = 116) and (hState = 582)) or
								((vState = 116) and (hState = 583)) or
								((vState = 116) and (hState = 584)) or
								((vState = 116) and (hState = 585)) or
								((vState = 116) and (hState = 586)) or
								((vState = 116) and (hState = 587)) or
								((vState = 116) and (hState = 592)) or
								((vState = 116) and (hState = 593)) or
								((vState = 116) and (hState = 594)) or
								((vState = 117) and (hState = 487)) or
								((vState = 117) and (hState = 488)) or
								((vState = 117) and (hState = 489)) or
								((vState = 117) and (hState = 490)) or
								((vState = 117) and (hState = 491)) or
								((vState = 117) and (hState = 492)) or
								((vState = 117) and (hState = 493)) or
								((vState = 117) and (hState = 494)) or
								((vState = 117) and (hState = 495)) or
								((vState = 117) and (hState = 496)) or
								((vState = 117) and (hState = 497)) or
								((vState = 117) and (hState = 498)) or
								((vState = 117) and (hState = 499)) or
								((vState = 117) and (hState = 500)) or
								((vState = 117) and (hState = 501)) or
								((vState = 117) and (hState = 502)) or
								((vState = 117) and (hState = 503)) or
								((vState = 117) and (hState = 505)) or
								((vState = 117) and (hState = 506)) or
								((vState = 117) and (hState = 507)) or
								((vState = 117) and (hState = 508)) or
								((vState = 117) and (hState = 509)) or
								((vState = 117) and (hState = 510)) or
								((vState = 117) and (hState = 511)) or
								((vState = 117) and (hState = 512)) or
								((vState = 117) and (hState = 513)) or
								((vState = 117) and (hState = 514)) or
								((vState = 117) and (hState = 516)) or
								((vState = 117) and (hState = 522)) or
								((vState = 117) and (hState = 523)) or
								((vState = 117) and (hState = 524)) or
								((vState = 117) and (hState = 525)) or
								((vState = 117) and (hState = 527)) or
								((vState = 117) and (hState = 528)) or
								((vState = 117) and (hState = 529)) or
								((vState = 117) and (hState = 534)) or
								((vState = 117) and (hState = 535)) or
								((vState = 117) and (hState = 536)) or
								((vState = 117) and (hState = 550)) or
								((vState = 117) and (hState = 551)) or
								((vState = 117) and (hState = 553)) or
								((vState = 117) and (hState = 554)) or
								((vState = 117) and (hState = 555)) or
								((vState = 117) and (hState = 559)) or
								((vState = 117) and (hState = 560)) or
								((vState = 117) and (hState = 561)) or
								((vState = 117) and (hState = 568)) or
								((vState = 117) and (hState = 569)) or
								((vState = 117) and (hState = 570)) or
								((vState = 117) and (hState = 575)) or
								((vState = 117) and (hState = 576)) or
								((vState = 117) and (hState = 577)) or
								((vState = 117) and (hState = 578)) or
								((vState = 117) and (hState = 581)) or
								((vState = 117) and (hState = 582)) or
								((vState = 117) and (hState = 583)) or
								((vState = 117) and (hState = 584)) or
								((vState = 117) and (hState = 585)) or
								((vState = 117) and (hState = 586)) or
								((vState = 117) and (hState = 591)) or
								((vState = 117) and (hState = 592)) or
								((vState = 117) and (hState = 593)) or
								((vState = 117) and (hState = 594)) or
								((vState = 118) and (hState = 488)) or
								((vState = 118) and (hState = 489)) or
								((vState = 118) and (hState = 490)) or
								((vState = 118) and (hState = 491)) or
								((vState = 118) and (hState = 492)) or
								((vState = 118) and (hState = 493)) or
								((vState = 118) and (hState = 505)) or
								((vState = 118) and (hState = 506)) or
								((vState = 118) and (hState = 507)) or
								((vState = 118) and (hState = 508)) or
								((vState = 118) and (hState = 509)) or
								((vState = 118) and (hState = 510)) or
								((vState = 118) and (hState = 511)) or
								((vState = 118) and (hState = 512)) or
								((vState = 118) and (hState = 513)) or
								((vState = 118) and (hState = 516)) or
								((vState = 118) and (hState = 520)) or
								((vState = 118) and (hState = 521)) or
								((vState = 118) and (hState = 522)) or
								((vState = 118) and (hState = 523)) or
								((vState = 118) and (hState = 526)) or
								((vState = 118) and (hState = 527)) or
								((vState = 118) and (hState = 528)) or
								((vState = 118) and (hState = 534)) or
								((vState = 118) and (hState = 535)) or
								((vState = 118) and (hState = 536)) or
								((vState = 118) and (hState = 537)) or
								((vState = 118) and (hState = 538)) or
								((vState = 118) and (hState = 550)) or
								((vState = 118) and (hState = 551)) or
								((vState = 118) and (hState = 552)) or
								((vState = 118) and (hState = 554)) or
								((vState = 118) and (hState = 555)) or
								((vState = 118) and (hState = 556)) or
								((vState = 118) and (hState = 557)) or
								((vState = 118) and (hState = 558)) or
								((vState = 118) and (hState = 559)) or
								((vState = 118) and (hState = 560)) or
								((vState = 118) and (hState = 561)) or
								((vState = 118) and (hState = 562)) or
								((vState = 118) and (hState = 563)) or
								((vState = 118) and (hState = 564)) or
								((vState = 118) and (hState = 565)) or
								((vState = 118) and (hState = 566)) or
								((vState = 118) and (hState = 567)) or
								((vState = 118) and (hState = 568)) or
								((vState = 118) and (hState = 569)) or
								((vState = 118) and (hState = 570)) or
								((vState = 118) and (hState = 571)) or
								((vState = 118) and (hState = 572)) or
								((vState = 118) and (hState = 573)) or
								((vState = 118) and (hState = 574)) or
								((vState = 118) and (hState = 575)) or
								((vState = 118) and (hState = 576)) or
								((vState = 118) and (hState = 577)) or
								((vState = 118) and (hState = 578)) or
								((vState = 118) and (hState = 579)) or
								((vState = 118) and (hState = 580)) or
								((vState = 118) and (hState = 581)) or
								((vState = 118) and (hState = 582)) or
								((vState = 118) and (hState = 583)) or
								((vState = 118) and (hState = 584)) or
								((vState = 118) and (hState = 585)) or
								((vState = 118) and (hState = 586)) or
								((vState = 118) and (hState = 591)) or
								((vState = 118) and (hState = 592)) or
								((vState = 118) and (hState = 593)) or
								((vState = 118) and (hState = 594)) or
								((vState = 118) and (hState = 598)) or
								((vState = 118) and (hState = 599)) or
								((vState = 119) and (hState = 489)) or
								((vState = 119) and (hState = 490)) or
								((vState = 119) and (hState = 492)) or
								((vState = 119) and (hState = 493)) or
								((vState = 119) and (hState = 494)) or
								((vState = 119) and (hState = 506)) or
								((vState = 119) and (hState = 507)) or
								((vState = 119) and (hState = 508)) or
								((vState = 119) and (hState = 509)) or
								((vState = 119) and (hState = 512)) or
								((vState = 119) and (hState = 513)) or
								((vState = 119) and (hState = 516)) or
								((vState = 119) and (hState = 518)) or
								((vState = 119) and (hState = 519)) or
								((vState = 119) and (hState = 520)) or
								((vState = 119) and (hState = 521)) or
								((vState = 119) and (hState = 522)) or
								((vState = 119) and (hState = 525)) or
								((vState = 119) and (hState = 526)) or
								((vState = 119) and (hState = 527)) or
								((vState = 119) and (hState = 534)) or
								((vState = 119) and (hState = 535)) or
								((vState = 119) and (hState = 536)) or
								((vState = 119) and (hState = 537)) or
								((vState = 119) and (hState = 538)) or
								((vState = 119) and (hState = 539)) or
								((vState = 119) and (hState = 540)) or
								((vState = 119) and (hState = 541)) or
								((vState = 119) and (hState = 551)) or
								((vState = 119) and (hState = 552)) or
								((vState = 119) and (hState = 553)) or
								((vState = 119) and (hState = 555)) or
								((vState = 119) and (hState = 556)) or
								((vState = 119) and (hState = 557)) or
								((vState = 119) and (hState = 558)) or
								((vState = 119) and (hState = 559)) or
								((vState = 119) and (hState = 560)) or
								((vState = 119) and (hState = 561)) or
								((vState = 119) and (hState = 562)) or
								((vState = 119) and (hState = 563)) or
								((vState = 119) and (hState = 564)) or
								((vState = 119) and (hState = 565)) or
								((vState = 119) and (hState = 566)) or
								((vState = 119) and (hState = 567)) or
								((vState = 119) and (hState = 568)) or
								((vState = 119) and (hState = 569)) or
								((vState = 119) and (hState = 570)) or
								((vState = 119) and (hState = 571)) or
								((vState = 119) and (hState = 572)) or
								((vState = 119) and (hState = 573)) or
								((vState = 119) and (hState = 574)) or
								((vState = 119) and (hState = 575)) or
								((vState = 119) and (hState = 576)) or
								((vState = 119) and (hState = 577)) or
								((vState = 119) and (hState = 578)) or
								((vState = 119) and (hState = 579)) or
								((vState = 119) and (hState = 580)) or
								((vState = 119) and (hState = 581)) or
								((vState = 119) and (hState = 582)) or
								((vState = 119) and (hState = 583)) or
								((vState = 119) and (hState = 584)) or
								((vState = 119) and (hState = 585)) or
								((vState = 119) and (hState = 586)) or
								((vState = 119) and (hState = 590)) or
								((vState = 119) and (hState = 591)) or
								((vState = 119) and (hState = 592)) or
								((vState = 119) and (hState = 593)) or
								((vState = 119) and (hState = 594)) or
								((vState = 119) and (hState = 598)) or
								((vState = 119) and (hState = 599)) or
								((vState = 120) and (hState = 490)) or
								((vState = 120) and (hState = 491)) or
								((vState = 120) and (hState = 493)) or
								((vState = 120) and (hState = 494)) or
								((vState = 120) and (hState = 495)) or
								((vState = 120) and (hState = 505)) or
								((vState = 120) and (hState = 506)) or
								((vState = 120) and (hState = 507)) or
								((vState = 120) and (hState = 508)) or
								((vState = 120) and (hState = 511)) or
								((vState = 120) and (hState = 512)) or
								((vState = 120) and (hState = 515)) or
								((vState = 120) and (hState = 516)) or
								((vState = 120) and (hState = 517)) or
								((vState = 120) and (hState = 518)) or
								((vState = 120) and (hState = 519)) or
								((vState = 120) and (hState = 520)) or
								((vState = 120) and (hState = 524)) or
								((vState = 120) and (hState = 525)) or
								((vState = 120) and (hState = 526)) or
								((vState = 120) and (hState = 537)) or
								((vState = 120) and (hState = 538)) or
								((vState = 120) and (hState = 539)) or
								((vState = 120) and (hState = 540)) or
								((vState = 120) and (hState = 541)) or
								((vState = 120) and (hState = 542)) or
								((vState = 120) and (hState = 543)) or
								((vState = 120) and (hState = 544)) or
								((vState = 120) and (hState = 545)) or
								((vState = 120) and (hState = 546)) or
								((vState = 120) and (hState = 547)) or
								((vState = 120) and (hState = 552)) or
								((vState = 120) and (hState = 553)) or
								((vState = 120) and (hState = 554)) or
								((vState = 120) and (hState = 555)) or
								((vState = 120) and (hState = 556)) or
								((vState = 120) and (hState = 557)) or
								((vState = 120) and (hState = 559)) or
								((vState = 120) and (hState = 560)) or
								((vState = 120) and (hState = 561)) or
								((vState = 120) and (hState = 562)) or
								((vState = 120) and (hState = 563)) or
								((vState = 120) and (hState = 564)) or
								((vState = 120) and (hState = 565)) or
								((vState = 120) and (hState = 566)) or
								((vState = 120) and (hState = 567)) or
								((vState = 120) and (hState = 568)) or
								((vState = 120) and (hState = 569)) or
								((vState = 120) and (hState = 570)) or
								((vState = 120) and (hState = 571)) or
								((vState = 120) and (hState = 572)) or
								((vState = 120) and (hState = 573)) or
								((vState = 120) and (hState = 574)) or
								((vState = 120) and (hState = 575)) or
								((vState = 120) and (hState = 576)) or
								((vState = 120) and (hState = 579)) or
								((vState = 120) and (hState = 580)) or
								((vState = 120) and (hState = 581)) or
								((vState = 120) and (hState = 582)) or
								((vState = 120) and (hState = 583)) or
								((vState = 120) and (hState = 584)) or
								((vState = 120) and (hState = 585)) or
								((vState = 120) and (hState = 586)) or
								((vState = 120) and (hState = 590)) or
								((vState = 120) and (hState = 591)) or
								((vState = 120) and (hState = 592)) or
								((vState = 120) and (hState = 593)) or
								((vState = 120) and (hState = 594)) or
								((vState = 120) and (hState = 596)) or
								((vState = 120) and (hState = 597)) or
								((vState = 120) and (hState = 598)) or
								((vState = 120) and (hState = 599)) or
								((vState = 121) and (hState = 490)) or
								((vState = 121) and (hState = 491)) or
								((vState = 121) and (hState = 492)) or
								((vState = 121) and (hState = 494)) or
								((vState = 121) and (hState = 495)) or
								((vState = 121) and (hState = 496)) or
								((vState = 121) and (hState = 504)) or
								((vState = 121) and (hState = 505)) or
								((vState = 121) and (hState = 506)) or
								((vState = 121) and (hState = 507)) or
								((vState = 121) and (hState = 508)) or
								((vState = 121) and (hState = 511)) or
								((vState = 121) and (hState = 512)) or
								((vState = 121) and (hState = 513)) or
								((vState = 121) and (hState = 514)) or
								((vState = 121) and (hState = 515)) or
								((vState = 121) and (hState = 516)) or
								((vState = 121) and (hState = 517)) or
								((vState = 121) and (hState = 518)) or
								((vState = 121) and (hState = 519)) or
								((vState = 121) and (hState = 520)) or
								((vState = 121) and (hState = 523)) or
								((vState = 121) and (hState = 524)) or
								((vState = 121) and (hState = 525)) or
								((vState = 121) and (hState = 539)) or
								((vState = 121) and (hState = 540)) or
								((vState = 121) and (hState = 541)) or
								((vState = 121) and (hState = 542)) or
								((vState = 121) and (hState = 543)) or
								((vState = 121) and (hState = 544)) or
								((vState = 121) and (hState = 545)) or
								((vState = 121) and (hState = 546)) or
								((vState = 121) and (hState = 547)) or
								((vState = 121) and (hState = 548)) or
								((vState = 121) and (hState = 549)) or
								((vState = 121) and (hState = 550)) or
								((vState = 121) and (hState = 551)) or
								((vState = 121) and (hState = 552)) or
								((vState = 121) and (hState = 553)) or
								((vState = 121) and (hState = 554)) or
								((vState = 121) and (hState = 555)) or
								((vState = 121) and (hState = 562)) or
								((vState = 121) and (hState = 563)) or
								((vState = 121) and (hState = 564)) or
								((vState = 121) and (hState = 565)) or
								((vState = 121) and (hState = 566)) or
								((vState = 121) and (hState = 567)) or
								((vState = 121) and (hState = 568)) or
								((vState = 121) and (hState = 569)) or
								((vState = 121) and (hState = 570)) or
								((vState = 121) and (hState = 571)) or
								((vState = 121) and (hState = 572)) or
								((vState = 121) and (hState = 573)) or
								((vState = 121) and (hState = 574)) or
								((vState = 121) and (hState = 575)) or
								((vState = 121) and (hState = 576)) or
								((vState = 121) and (hState = 577)) or
								((vState = 121) and (hState = 578)) or
								((vState = 121) and (hState = 579)) or
								((vState = 121) and (hState = 580)) or
								((vState = 121) and (hState = 584)) or
								((vState = 121) and (hState = 585)) or
								((vState = 121) and (hState = 586)) or
								((vState = 121) and (hState = 587)) or
								((vState = 121) and (hState = 588)) or
								((vState = 121) and (hState = 589)) or
								((vState = 121) and (hState = 590)) or
								((vState = 121) and (hState = 591)) or
								((vState = 121) and (hState = 592)) or
								((vState = 121) and (hState = 593)) or
								((vState = 121) and (hState = 594)) or
								((vState = 121) and (hState = 595)) or
								((vState = 121) and (hState = 596)) or
								((vState = 121) and (hState = 597)) or
								((vState = 121) and (hState = 598)) or
								((vState = 122) and (hState = 491)) or
								((vState = 122) and (hState = 492)) or
								((vState = 122) and (hState = 495)) or
								((vState = 122) and (hState = 496)) or
								((vState = 122) and (hState = 497)) or
								((vState = 122) and (hState = 502)) or
								((vState = 122) and (hState = 503)) or
								((vState = 122) and (hState = 504)) or
								((vState = 122) and (hState = 505)) or
								((vState = 122) and (hState = 508)) or
								((vState = 122) and (hState = 509)) or
								((vState = 122) and (hState = 510)) or
								((vState = 122) and (hState = 511)) or
								((vState = 122) and (hState = 512)) or
								((vState = 122) and (hState = 513)) or
								((vState = 122) and (hState = 514)) or
								((vState = 122) and (hState = 515)) or
								((vState = 122) and (hState = 516)) or
								((vState = 122) and (hState = 517)) or
								((vState = 122) and (hState = 518)) or
								((vState = 122) and (hState = 519)) or
								((vState = 122) and (hState = 520)) or
								((vState = 122) and (hState = 523)) or
								((vState = 122) and (hState = 524)) or
								((vState = 122) and (hState = 541)) or
								((vState = 122) and (hState = 542)) or
								((vState = 122) and (hState = 543)) or
								((vState = 122) and (hState = 548)) or
								((vState = 122) and (hState = 549)) or
								((vState = 122) and (hState = 550)) or
								((vState = 122) and (hState = 551)) or
								((vState = 122) and (hState = 552)) or
								((vState = 122) and (hState = 553)) or
								((vState = 122) and (hState = 554)) or
								((vState = 122) and (hState = 555)) or
								((vState = 122) and (hState = 561)) or
								((vState = 122) and (hState = 562)) or
								((vState = 122) and (hState = 563)) or
								((vState = 122) and (hState = 567)) or
								((vState = 122) and (hState = 568)) or
								((vState = 122) and (hState = 569)) or
								((vState = 122) and (hState = 570)) or
								((vState = 122) and (hState = 572)) or
								((vState = 122) and (hState = 573)) or
								((vState = 122) and (hState = 574)) or
								((vState = 122) and (hState = 575)) or
								((vState = 122) and (hState = 576)) or
								((vState = 122) and (hState = 577)) or
								((vState = 122) and (hState = 578)) or
								((vState = 122) and (hState = 579)) or
								((vState = 122) and (hState = 580)) or
								((vState = 122) and (hState = 581)) or
								((vState = 122) and (hState = 582)) or
								((vState = 122) and (hState = 583)) or
								((vState = 122) and (hState = 584)) or
								((vState = 122) and (hState = 585)) or
								((vState = 122) and (hState = 586)) or
								((vState = 122) and (hState = 587)) or
								((vState = 122) and (hState = 588)) or
								((vState = 122) and (hState = 589)) or
								((vState = 122) and (hState = 590)) or
								((vState = 122) and (hState = 591)) or
								((vState = 122) and (hState = 592)) or
								((vState = 122) and (hState = 593)) or
								((vState = 122) and (hState = 594)) or
								((vState = 122) and (hState = 595)) or
								((vState = 122) and (hState = 596)) or
								((vState = 122) and (hState = 597)) or
								((vState = 122) and (hState = 598)) or
								((vState = 123) and (hState = 492)) or
								((vState = 123) and (hState = 493)) or
								((vState = 123) and (hState = 496)) or
								((vState = 123) and (hState = 497)) or
								((vState = 123) and (hState = 498)) or
								((vState = 123) and (hState = 500)) or
								((vState = 123) and (hState = 501)) or
								((vState = 123) and (hState = 502)) or
								((vState = 123) and (hState = 503)) or
								((vState = 123) and (hState = 509)) or
								((vState = 123) and (hState = 510)) or
								((vState = 123) and (hState = 511)) or
								((vState = 123) and (hState = 512)) or
								((vState = 123) and (hState = 513)) or
								((vState = 123) and (hState = 514)) or
								((vState = 123) and (hState = 516)) or
								((vState = 123) and (hState = 517)) or
								((vState = 123) and (hState = 518)) or
								((vState = 123) and (hState = 519)) or
								((vState = 123) and (hState = 522)) or
								((vState = 123) and (hState = 523)) or
								((vState = 123) and (hState = 542)) or
								((vState = 123) and (hState = 543)) or
								((vState = 123) and (hState = 544)) or
								((vState = 123) and (hState = 545)) or
								((vState = 123) and (hState = 552)) or
								((vState = 123) and (hState = 555)) or
								((vState = 123) and (hState = 556)) or
								((vState = 123) and (hState = 559)) or
								((vState = 123) and (hState = 560)) or
								((vState = 123) and (hState = 561)) or
								((vState = 123) and (hState = 562)) or
								((vState = 123) and (hState = 565)) or
								((vState = 123) and (hState = 566)) or
								((vState = 123) and (hState = 567)) or
								((vState = 123) and (hState = 568)) or
								((vState = 123) and (hState = 574)) or
								((vState = 123) and (hState = 575)) or
								((vState = 123) and (hState = 576)) or
								((vState = 123) and (hState = 577)) or
								((vState = 123) and (hState = 578)) or
								((vState = 123) and (hState = 579)) or
								((vState = 123) and (hState = 580)) or
								((vState = 123) and (hState = 581)) or
								((vState = 123) and (hState = 582)) or
								((vState = 123) and (hState = 583)) or
								((vState = 123) and (hState = 584)) or
								((vState = 123) and (hState = 585)) or
								((vState = 123) and (hState = 586)) or
								((vState = 123) and (hState = 587)) or
								((vState = 123) and (hState = 588)) or
								((vState = 123) and (hState = 589)) or
								((vState = 123) and (hState = 590)) or
								((vState = 123) and (hState = 591)) or
								((vState = 123) and (hState = 592)) or
								((vState = 123) and (hState = 593)) or
								((vState = 123) and (hState = 594)) or
								((vState = 123) and (hState = 595)) or
								((vState = 123) and (hState = 596)) or
								((vState = 123) and (hState = 597)) or
								((vState = 124) and (hState = 493)) or
								((vState = 124) and (hState = 494)) or
								((vState = 124) and (hState = 495)) or
								((vState = 124) and (hState = 497)) or
								((vState = 124) and (hState = 498)) or
								((vState = 124) and (hState = 499)) or
								((vState = 124) and (hState = 500)) or
								((vState = 124) and (hState = 501)) or
								((vState = 124) and (hState = 509)) or
								((vState = 124) and (hState = 510)) or
								((vState = 124) and (hState = 511)) or
								((vState = 124) and (hState = 515)) or
								((vState = 124) and (hState = 516)) or
								((vState = 124) and (hState = 517)) or
								((vState = 124) and (hState = 520)) or
								((vState = 124) and (hState = 521)) or
								((vState = 124) and (hState = 522)) or
								((vState = 124) and (hState = 545)) or
								((vState = 124) and (hState = 546)) or
								((vState = 124) and (hState = 547)) or
								((vState = 124) and (hState = 556)) or
								((vState = 124) and (hState = 557)) or
								((vState = 124) and (hState = 558)) or
								((vState = 124) and (hState = 559)) or
								((vState = 124) and (hState = 560)) or
								((vState = 124) and (hState = 564)) or
								((vState = 124) and (hState = 565)) or
								((vState = 124) and (hState = 566)) or
								((vState = 124) and (hState = 574)) or
								((vState = 124) and (hState = 575)) or
								((vState = 124) and (hState = 576)) or
								((vState = 124) and (hState = 577)) or
								((vState = 124) and (hState = 578)) or
								((vState = 124) and (hState = 587)) or
								((vState = 124) and (hState = 588)) or
								((vState = 124) and (hState = 589)) or
								((vState = 124) and (hState = 590)) or
								((vState = 124) and (hState = 591)) or
								((vState = 124) and (hState = 592)) or
								((vState = 124) and (hState = 593)) or
								((vState = 124) and (hState = 594)) or
								((vState = 124) and (hState = 595)) or
								((vState = 125) and (hState = 493)) or
								((vState = 125) and (hState = 494)) or
								((vState = 125) and (hState = 495)) or
								((vState = 125) and (hState = 496)) or
								((vState = 125) and (hState = 497)) or
								((vState = 125) and (hState = 498)) or
								((vState = 125) and (hState = 499)) or
								((vState = 125) and (hState = 500)) or
								((vState = 125) and (hState = 501)) or
								((vState = 125) and (hState = 507)) or
								((vState = 125) and (hState = 508)) or
								((vState = 125) and (hState = 509)) or
								((vState = 125) and (hState = 510)) or
								((vState = 125) and (hState = 511)) or
								((vState = 125) and (hState = 514)) or
								((vState = 125) and (hState = 515)) or
								((vState = 125) and (hState = 516)) or
								((vState = 125) and (hState = 517)) or
								((vState = 125) and (hState = 519)) or
								((vState = 125) and (hState = 520)) or
								((vState = 125) and (hState = 521)) or
								((vState = 125) and (hState = 546)) or
								((vState = 125) and (hState = 547)) or
								((vState = 125) and (hState = 548)) or
								((vState = 125) and (hState = 549)) or
								((vState = 125) and (hState = 556)) or
								((vState = 125) and (hState = 557)) or
								((vState = 125) and (hState = 558)) or
								((vState = 125) and (hState = 559)) or
								((vState = 125) and (hState = 560)) or
								((vState = 125) and (hState = 563)) or
								((vState = 125) and (hState = 564)) or
								((vState = 125) and (hState = 565)) or
								((vState = 125) and (hState = 566)) or
								((vState = 125) and (hState = 574)) or
								((vState = 125) and (hState = 575)) or
								((vState = 125) and (hState = 576)) or
								((vState = 125) and (hState = 577)) or
								((vState = 125) and (hState = 587)) or
								((vState = 125) and (hState = 588)) or
								((vState = 125) and (hState = 590)) or
								((vState = 125) and (hState = 591)) or
								((vState = 125) and (hState = 592)) or
								((vState = 125) and (hState = 593)) or
								((vState = 125) and (hState = 594)) or
								((vState = 125) and (hState = 595)) or
								((vState = 125) and (hState = 596)) or
								((vState = 126) and (hState = 496)) or
								((vState = 126) and (hState = 497)) or
								((vState = 126) and (hState = 498)) or
								((vState = 126) and (hState = 499)) or
								((vState = 126) and (hState = 500)) or
								((vState = 126) and (hState = 501)) or
								((vState = 126) and (hState = 502)) or
								((vState = 126) and (hState = 503)) or
								((vState = 126) and (hState = 504)) or
								((vState = 126) and (hState = 505)) or
								((vState = 126) and (hState = 506)) or
								((vState = 126) and (hState = 507)) or
								((vState = 126) and (hState = 508)) or
								((vState = 126) and (hState = 510)) or
								((vState = 126) and (hState = 511)) or
								((vState = 126) and (hState = 512)) or
								((vState = 126) and (hState = 513)) or
								((vState = 126) and (hState = 514)) or
								((vState = 126) and (hState = 515)) or
								((vState = 126) and (hState = 516)) or
								((vState = 126) and (hState = 517)) or
								((vState = 126) and (hState = 518)) or
								((vState = 126) and (hState = 519)) or
								((vState = 126) and (hState = 520)) or
								((vState = 126) and (hState = 548)) or
								((vState = 126) and (hState = 549)) or
								((vState = 126) and (hState = 550)) or
								((vState = 126) and (hState = 551)) or
								((vState = 126) and (hState = 557)) or
								((vState = 126) and (hState = 558)) or
								((vState = 126) and (hState = 559)) or
								((vState = 126) and (hState = 560)) or
								((vState = 126) and (hState = 561)) or
								((vState = 126) and (hState = 563)) or
								((vState = 126) and (hState = 564)) or
								((vState = 126) and (hState = 565)) or
								((vState = 126) and (hState = 566)) or
								((vState = 126) and (hState = 567)) or
								((vState = 126) and (hState = 568)) or
								((vState = 126) and (hState = 569)) or
								((vState = 126) and (hState = 570)) or
								((vState = 126) and (hState = 571)) or
								((vState = 126) and (hState = 573)) or
								((vState = 126) and (hState = 574)) or
								((vState = 126) and (hState = 575)) or
								((vState = 126) and (hState = 576)) or
								((vState = 126) and (hState = 577)) or
								((vState = 126) and (hState = 586)) or
								((vState = 126) and (hState = 587)) or
								((vState = 126) and (hState = 588)) or
								((vState = 126) and (hState = 589)) or
								((vState = 126) and (hState = 590)) or
								((vState = 126) and (hState = 591)) or
								((vState = 126) and (hState = 592)) or
								((vState = 126) and (hState = 595)) or
								((vState = 126) and (hState = 596)) or
								((vState = 126) and (hState = 597)) or
								((vState = 126) and (hState = 598)) or
								((vState = 127) and (hState = 505)) or
								((vState = 127) and (hState = 506)) or
								((vState = 127) and (hState = 511)) or
								((vState = 127) and (hState = 512)) or
								((vState = 127) and (hState = 513)) or
								((vState = 127) and (hState = 516)) or
								((vState = 127) and (hState = 517)) or
								((vState = 127) and (hState = 518)) or
								((vState = 127) and (hState = 519)) or
								((vState = 127) and (hState = 550)) or
								((vState = 127) and (hState = 551)) or
								((vState = 127) and (hState = 552)) or
								((vState = 127) and (hState = 553)) or
								((vState = 127) and (hState = 558)) or
								((vState = 127) and (hState = 559)) or
								((vState = 127) and (hState = 560)) or
								((vState = 127) and (hState = 561)) or
								((vState = 127) and (hState = 562)) or
								((vState = 127) and (hState = 563)) or
								((vState = 127) and (hState = 567)) or
								((vState = 127) and (hState = 568)) or
								((vState = 127) and (hState = 569)) or
								((vState = 127) and (hState = 570)) or
								((vState = 127) and (hState = 571)) or
								((vState = 127) and (hState = 572)) or
								((vState = 127) and (hState = 573)) or
								((vState = 127) and (hState = 574)) or
								((vState = 127) and (hState = 575)) or
								((vState = 127) and (hState = 576)) or
								((vState = 127) and (hState = 577)) or
								((vState = 127) and (hState = 578)) or
								((vState = 127) and (hState = 579)) or
								((vState = 127) and (hState = 586)) or
								((vState = 127) and (hState = 587)) or
								((vState = 127) and (hState = 588)) or
								((vState = 127) and (hState = 589)) or
								((vState = 127) and (hState = 590)) or
								((vState = 127) and (hState = 591)) or
								((vState = 127) and (hState = 592)) or
								((vState = 127) and (hState = 595)) or
								((vState = 127) and (hState = 596)) or
								((vState = 127) and (hState = 597)) or
								((vState = 127) and (hState = 598)) or
								((vState = 127) and (hState = 599)) or
								((vState = 128) and (hState = 516)) or
								((vState = 128) and (hState = 517)) or
								((vState = 128) and (hState = 518)) or
								((vState = 128) and (hState = 552)) or
								((vState = 128) and (hState = 553)) or
								((vState = 128) and (hState = 554)) or
								((vState = 128) and (hState = 559)) or
								((vState = 128) and (hState = 560)) or
								((vState = 128) and (hState = 562)) or
								((vState = 128) and (hState = 563)) or
								((vState = 128) and (hState = 564)) or
								((vState = 128) and (hState = 568)) or
								((vState = 128) and (hState = 569)) or
								((vState = 128) and (hState = 570)) or
								((vState = 128) and (hState = 571)) or
								((vState = 128) and (hState = 572)) or
								((vState = 128) and (hState = 573)) or
								((vState = 128) and (hState = 574)) or
								((vState = 128) and (hState = 575)) or
								((vState = 128) and (hState = 576)) or
								((vState = 128) and (hState = 577)) or
								((vState = 128) and (hState = 578)) or
								((vState = 128) and (hState = 579)) or
								((vState = 128) and (hState = 580)) or
								((vState = 128) and (hState = 585)) or
								((vState = 128) and (hState = 586)) or
								((vState = 128) and (hState = 587)) or
								((vState = 128) and (hState = 588)) or
								((vState = 128) and (hState = 589)) or
								((vState = 128) and (hState = 590)) or
								((vState = 128) and (hState = 591)) or
								((vState = 128) and (hState = 592)) or
								((vState = 128) and (hState = 593)) or
								((vState = 128) and (hState = 594)) or
								((vState = 128) and (hState = 595)) or
								((vState = 128) and (hState = 596)) or
								((vState = 128) and (hState = 597)) or
								((vState = 128) and (hState = 598)) or
								((vState = 129) and (hState = 517)) or
								((vState = 129) and (hState = 553)) or
								((vState = 129) and (hState = 554)) or
								((vState = 129) and (hState = 555)) or
								((vState = 129) and (hState = 556)) or
								((vState = 129) and (hState = 560)) or
								((vState = 129) and (hState = 561)) or
								((vState = 129) and (hState = 563)) or
								((vState = 129) and (hState = 564)) or
								((vState = 129) and (hState = 565)) or
								((vState = 129) and (hState = 572)) or
								((vState = 129) and (hState = 573)) or
								((vState = 129) and (hState = 574)) or
								((vState = 129) and (hState = 577)) or
								((vState = 129) and (hState = 578)) or
								((vState = 129) and (hState = 579)) or
								((vState = 129) and (hState = 584)) or
								((vState = 129) and (hState = 585)) or
								((vState = 129) and (hState = 586)) or
								((vState = 129) and (hState = 587)) or
								((vState = 129) and (hState = 588)) or
								((vState = 129) and (hState = 589)) or
								((vState = 129) and (hState = 590)) or
								((vState = 129) and (hState = 591)) or
								((vState = 129) and (hState = 592)) or
								((vState = 129) and (hState = 593)) or
								((vState = 129) and (hState = 594)) or
								((vState = 130) and (hState = 555)) or
								((vState = 130) and (hState = 556)) or
								((vState = 130) and (hState = 557)) or
								((vState = 130) and (hState = 560)) or
								((vState = 130) and (hState = 561)) or
								((vState = 130) and (hState = 564)) or
								((vState = 130) and (hState = 565)) or
								((vState = 130) and (hState = 566)) or
								((vState = 130) and (hState = 572)) or
								((vState = 130) and (hState = 573)) or
								((vState = 130) and (hState = 584)) or
								((vState = 130) and (hState = 585)) or
								((vState = 130) and (hState = 586)) or
								((vState = 130) and (hState = 587)) or
								((vState = 130) and (hState = 588)) or
								((vState = 130) and (hState = 590)) or
								((vState = 130) and (hState = 591)) or
								((vState = 131) and (hState = 556)) or
								((vState = 131) and (hState = 557)) or
								((vState = 131) and (hState = 561)) or
								((vState = 131) and (hState = 562)) or
								((vState = 131) and (hState = 566)) or
								((vState = 131) and (hState = 567)) or
								((vState = 131) and (hState = 572)) or
								((vState = 131) and (hState = 573)) or
								((vState = 131) and (hState = 584)) or
								((vState = 131) and (hState = 585)) or
								((vState = 131) and (hState = 586)) or
								((vState = 131) and (hState = 587)) or
								((vState = 131) and (hState = 590)) or
								((vState = 131) and (hState = 591)) or
								((vState = 132) and (hState = 556)) or
								((vState = 132) and (hState = 557)) or
								((vState = 132) and (hState = 561)) or
								((vState = 132) and (hState = 562)) or
								((vState = 132) and (hState = 567)) or
								((vState = 132) and (hState = 568)) or
								((vState = 132) and (hState = 569)) or
								((vState = 132) and (hState = 572)) or
								((vState = 132) and (hState = 583)) or
								((vState = 132) and (hState = 584)) or
								((vState = 132) and (hState = 585)) or
								((vState = 132) and (hState = 586)) or
								((vState = 132) and (hState = 597)) or
								((vState = 133) and (hState = 557)) or
								((vState = 133) and (hState = 558)) or
								((vState = 133) and (hState = 562)) or
								((vState = 133) and (hState = 563)) or
								((vState = 133) and (hState = 568)) or
								((vState = 133) and (hState = 569)) or
								((vState = 133) and (hState = 570)) or
								((vState = 133) and (hState = 571)) or
								((vState = 133) and (hState = 572)) or
								((vState = 133) and (hState = 583)) or
								((vState = 133) and (hState = 584)) or
								((vState = 133) and (hState = 585)) or
								((vState = 133) and (hState = 586)) or
								((vState = 133) and (hState = 590)) or
								((vState = 133) and (hState = 591)) or
								((vState = 133) and (hState = 592)) or
								((vState = 133) and (hState = 593)) or
								((vState = 133) and (hState = 594)) or
								((vState = 133) and (hState = 595)) or
								((vState = 133) and (hState = 596)) or
								((vState = 133) and (hState = 597)) or
								((vState = 133) and (hState = 598)) or
								((vState = 134) and (hState = 557)) or
								((vState = 134) and (hState = 558)) or
								((vState = 134) and (hState = 562)) or
								((vState = 134) and (hState = 563)) or
								((vState = 134) and (hState = 569)) or
								((vState = 134) and (hState = 570)) or
								((vState = 134) and (hState = 571)) or
								((vState = 134) and (hState = 572)) or
								((vState = 134) and (hState = 573)) or
								((vState = 134) and (hState = 582)) or
								((vState = 134) and (hState = 583)) or
								((vState = 134) and (hState = 584)) or
								((vState = 134) and (hState = 585)) or
								((vState = 134) and (hState = 586)) or
								((vState = 134) and (hState = 587)) or
								((vState = 134) and (hState = 588)) or
								((vState = 134) and (hState = 589)) or
								((vState = 134) and (hState = 590)) or
								((vState = 134) and (hState = 591)) or
								((vState = 134) and (hState = 592)) or
								((vState = 134) and (hState = 593)) or
								((vState = 134) and (hState = 596)) or
								((vState = 134) and (hState = 597)) or
								((vState = 134) and (hState = 598)) or
								((vState = 135) and (hState = 557)) or
								((vState = 135) and (hState = 558)) or
								((vState = 135) and (hState = 562)) or
								((vState = 135) and (hState = 563)) or
								((vState = 135) and (hState = 570)) or
								((vState = 135) and (hState = 571)) or
								((vState = 135) and (hState = 572)) or
								((vState = 135) and (hState = 573)) or
								((vState = 135) and (hState = 574)) or
								((vState = 135) and (hState = 578)) or
								((vState = 135) and (hState = 579)) or
								((vState = 135) and (hState = 580)) or
								((vState = 135) and (hState = 581)) or
								((vState = 135) and (hState = 582)) or
								((vState = 135) and (hState = 583)) or
								((vState = 135) and (hState = 584)) or
								((vState = 135) and (hState = 585)) or
								((vState = 135) and (hState = 586)) or
								((vState = 135) and (hState = 587)) or
								((vState = 135) and (hState = 588)) or
								((vState = 135) and (hState = 589)) or
								((vState = 135) and (hState = 596)) or
								((vState = 135) and (hState = 597)) or
								((vState = 136) and (hState = 557)) or
								((vState = 136) and (hState = 558)) or
								((vState = 136) and (hState = 562)) or
								((vState = 136) and (hState = 563)) or
								((vState = 136) and (hState = 572)) or
								((vState = 136) and (hState = 573)) or
								((vState = 136) and (hState = 574)) or
								((vState = 136) and (hState = 575)) or
								((vState = 136) and (hState = 576)) or
								((vState = 136) and (hState = 577)) or
								((vState = 136) and (hState = 578)) or
								((vState = 136) and (hState = 579)) or
								((vState = 136) and (hState = 580)) or
								((vState = 136) and (hState = 581)) or
								((vState = 136) and (hState = 582)) or
								((vState = 136) and (hState = 583)) or
								((vState = 136) and (hState = 596)) or
								((vState = 136) and (hState = 597)) or
								((vState = 137) and (hState = 558)) or
								((vState = 137) and (hState = 559)) or
								((vState = 137) and (hState = 563)) or
								((vState = 137) and (hState = 564)) or
								((vState = 137) and (hState = 573)) or
								((vState = 137) and (hState = 574)) or
								((vState = 137) and (hState = 575)) or
								((vState = 137) and (hState = 576)) or
								((vState = 137) and (hState = 577)) or
								((vState = 137) and (hState = 578)) or
								((vState = 137) and (hState = 581)) or
								((vState = 137) and (hState = 585)) or
								((vState = 137) and (hState = 586)) or
								((vState = 137) and (hState = 587)) or
								((vState = 137) and (hState = 596)) or
								((vState = 138) and (hState = 558)) or
								((vState = 138) and (hState = 559)) or
								((vState = 138) and (hState = 563)) or
								((vState = 138) and (hState = 564)) or
								((vState = 138) and (hState = 574)) or
								((vState = 138) and (hState = 575)) or
								((vState = 138) and (hState = 576)) or
								((vState = 138) and (hState = 577)) or
								((vState = 138) and (hState = 578)) or
								((vState = 138) and (hState = 584)) or
								((vState = 138) and (hState = 585)) or
								((vState = 138) and (hState = 586)) or
								((vState = 138) and (hState = 587)) or
								((vState = 138) and (hState = 595)) or
								((vState = 138) and (hState = 596)) or
								((vState = 138) and (hState = 599)) or
								((vState = 139) and (hState = 559)) or
								((vState = 139) and (hState = 563)) or
								((vState = 139) and (hState = 564)) or
								((vState = 139) and (hState = 572)) or
								((vState = 139) and (hState = 576)) or
								((vState = 139) and (hState = 577)) or
								((vState = 139) and (hState = 578)) or
								((vState = 139) and (hState = 579)) or
								((vState = 139) and (hState = 582)) or
								((vState = 139) and (hState = 583)) or
								((vState = 139) and (hState = 584)) or
								((vState = 139) and (hState = 585)) or
								((vState = 139) and (hState = 586)) or
								((vState = 139) and (hState = 590)) or
								((vState = 139) and (hState = 591)) or
								((vState = 139) and (hState = 592)) or
								((vState = 139) and (hState = 595)) or
								((vState = 139) and (hState = 596)) or
								((vState = 139) and (hState = 597)) or
								((vState = 139) and (hState = 598)) or
								((vState = 139) and (hState = 599)) or
								((vState = 140) and (hState = 559)) or
								((vState = 140) and (hState = 560)) or
								((vState = 140) and (hState = 564)) or
								((vState = 140) and (hState = 571)) or
								((vState = 140) and (hState = 572)) or
								((vState = 140) and (hState = 577)) or
								((vState = 140) and (hState = 578)) or
								((vState = 140) and (hState = 579)) or
								((vState = 140) and (hState = 580)) or
								((vState = 140) and (hState = 581)) or
								((vState = 140) and (hState = 582)) or
								((vState = 140) and (hState = 583)) or
								((vState = 140) and (hState = 584)) or
								((vState = 140) and (hState = 589)) or
								((vState = 140) and (hState = 590)) or
								((vState = 140) and (hState = 591)) or
								((vState = 140) and (hState = 592)) or
								((vState = 140) and (hState = 595)) or
								((vState = 140) and (hState = 596)) or
								((vState = 140) and (hState = 597)) or
								((vState = 140) and (hState = 598)) or
								((vState = 140) and (hState = 599)) or
								((vState = 141) and (hState = 559)) or
								((vState = 141) and (hState = 560)) or
								((vState = 141) and (hState = 564)) or
								((vState = 141) and (hState = 565)) or
								((vState = 141) and (hState = 570)) or
								((vState = 141) and (hState = 571)) or
								((vState = 141) and (hState = 572)) or
								((vState = 141) and (hState = 578)) or
								((vState = 141) and (hState = 579)) or
								((vState = 141) and (hState = 580)) or
								((vState = 141) and (hState = 581)) or
								((vState = 141) and (hState = 582)) or
								((vState = 141) and (hState = 583)) or
								((vState = 141) and (hState = 587)) or
								((vState = 141) and (hState = 588)) or
								((vState = 141) and (hState = 589)) or
								((vState = 141) and (hState = 590)) or
								((vState = 141) and (hState = 591)) or
								((vState = 141) and (hState = 594)) or
								((vState = 141) and (hState = 595)) or
								((vState = 141) and (hState = 596)) or
								((vState = 141) and (hState = 597)) or
								((vState = 141) and (hState = 599)) or
								((vState = 142) and (hState = 559)) or
								((vState = 142) and (hState = 560)) or
								((vState = 142) and (hState = 564)) or
								((vState = 142) and (hState = 565)) or
								((vState = 142) and (hState = 569)) or
								((vState = 142) and (hState = 570)) or
								((vState = 142) and (hState = 571)) or
								((vState = 142) and (hState = 572)) or
								((vState = 142) and (hState = 576)) or
								((vState = 142) and (hState = 577)) or
								((vState = 142) and (hState = 578)) or
								((vState = 142) and (hState = 579)) or
								((vState = 142) and (hState = 580)) or
								((vState = 142) and (hState = 581)) or
								((vState = 142) and (hState = 582)) or
								((vState = 142) and (hState = 586)) or
								((vState = 142) and (hState = 587)) or
								((vState = 142) and (hState = 588)) or
								((vState = 142) and (hState = 589)) or
								((vState = 142) and (hState = 590)) or
								((vState = 142) and (hState = 594)) or
								((vState = 142) and (hState = 595)) or
								((vState = 142) and (hState = 596)) or
								((vState = 142) and (hState = 597)) or
								((vState = 142) and (hState = 599)) or
								((vState = 143) and (hState = 560)) or
								((vState = 143) and (hState = 561)) or
								((vState = 143) and (hState = 564)) or
								((vState = 143) and (hState = 565)) or
								((vState = 143) and (hState = 569)) or
								((vState = 143) and (hState = 570)) or
								((vState = 143) and (hState = 572)) or
								((vState = 143) and (hState = 573)) or
								((vState = 143) and (hState = 574)) or
								((vState = 143) and (hState = 575)) or
								((vState = 143) and (hState = 576)) or
								((vState = 143) and (hState = 577)) or
								((vState = 143) and (hState = 578)) or
								((vState = 143) and (hState = 579)) or
								((vState = 143) and (hState = 580)) or
								((vState = 143) and (hState = 581)) or
								((vState = 143) and (hState = 582)) or
								((vState = 143) and (hState = 583)) or
								((vState = 143) and (hState = 584)) or
								((vState = 143) and (hState = 585)) or
								((vState = 143) and (hState = 586)) or
								((vState = 143) and (hState = 587)) or
								((vState = 143) and (hState = 588)) or
								((vState = 143) and (hState = 589)) or
								((vState = 143) and (hState = 590)) or
								((vState = 143) and (hState = 592)) or
								((vState = 143) and (hState = 593)) or
								((vState = 143) and (hState = 594)) or
								((vState = 143) and (hState = 595)) or
								((vState = 143) and (hState = 596)) or
								((vState = 143) and (hState = 599)) or
								((vState = 144) and (hState = 560)) or
								((vState = 144) and (hState = 561)) or
								((vState = 144) and (hState = 562)) or
								((vState = 144) and (hState = 563)) or
								((vState = 144) and (hState = 564)) or
								((vState = 144) and (hState = 565)) or
								((vState = 144) and (hState = 566)) or
								((vState = 144) and (hState = 567)) or
								((vState = 144) and (hState = 568)) or
								((vState = 144) and (hState = 569)) or
								((vState = 144) and (hState = 570)) or
								((vState = 144) and (hState = 571)) or
								((vState = 144) and (hState = 572)) or
								((vState = 144) and (hState = 573)) or
								((vState = 144) and (hState = 574)) or
								((vState = 144) and (hState = 575)) or
								((vState = 144) and (hState = 576)) or
								((vState = 144) and (hState = 577)) or
								((vState = 144) and (hState = 578)) or
								((vState = 144) and (hState = 579)) or
								((vState = 144) and (hState = 580)) or
								((vState = 144) and (hState = 581)) or
								((vState = 144) and (hState = 582)) or
								((vState = 144) and (hState = 583)) or
								((vState = 144) and (hState = 584)) or
								((vState = 144) and (hState = 585)) or
								((vState = 144) and (hState = 586)) or
								((vState = 144) and (hState = 587)) or
								((vState = 144) and (hState = 588)) or
								((vState = 144) and (hState = 589)) or
								((vState = 144) and (hState = 590)) or
								((vState = 144) and (hState = 591)) or
								((vState = 144) and (hState = 592)) or
								((vState = 144) and (hState = 593)) or
								((vState = 144) and (hState = 594)) or
								((vState = 144) and (hState = 595)) or
								((vState = 144) and (hState = 597)) or
								((vState = 144) and (hState = 599)) or
								((vState = 145) and (hState = 555)) or
								((vState = 145) and (hState = 556)) or
								((vState = 145) and (hState = 557)) or
								((vState = 145) and (hState = 558)) or
								((vState = 145) and (hState = 559)) or
								((vState = 145) and (hState = 560)) or
								((vState = 145) and (hState = 561)) or
								((vState = 145) and (hState = 562)) or
								((vState = 145) and (hState = 563)) or
								((vState = 145) and (hState = 564)) or
								((vState = 145) and (hState = 565)) or
								((vState = 145) and (hState = 566)) or
								((vState = 145) and (hState = 567)) or
								((vState = 145) and (hState = 568)) or
								((vState = 145) and (hState = 569)) or
								((vState = 145) and (hState = 570)) or
								((vState = 145) and (hState = 571)) or
								((vState = 145) and (hState = 572)) or
								((vState = 145) and (hState = 573)) or
								((vState = 145) and (hState = 574)) or
								((vState = 145) and (hState = 575)) or
								((vState = 145) and (hState = 576)) or
								((vState = 145) and (hState = 577)) or
								((vState = 145) and (hState = 578)) or
								((vState = 145) and (hState = 579)) or
								((vState = 145) and (hState = 580)) or
								((vState = 145) and (hState = 581)) or
								((vState = 145) and (hState = 582)) or
								((vState = 145) and (hState = 583)) or
								((vState = 145) and (hState = 584)) or
								((vState = 145) and (hState = 585)) or
								((vState = 145) and (hState = 586)) or
								((vState = 145) and (hState = 587)) or
								((vState = 145) and (hState = 588)) or
								((vState = 145) and (hState = 589)) or
								((vState = 145) and (hState = 590)) or
								((vState = 145) and (hState = 591)) or
								((vState = 145) and (hState = 592)) or
								((vState = 145) and (hState = 593)) or
								((vState = 145) and (hState = 594)) or
								((vState = 145) and (hState = 595)) or
								((vState = 145) and (hState = 596)) or
								((vState = 145) and (hState = 597)) or
								((vState = 145) and (hState = 598)) or
								((vState = 145) and (hState = 599)) or
								((vState = 146) and (hState = 555)) or
								((vState = 146) and (hState = 556)) or
								((vState = 146) and (hState = 557)) or
								((vState = 146) and (hState = 558)) or
								((vState = 146) and (hState = 559)) or
								((vState = 146) and (hState = 560)) or
								((vState = 146) and (hState = 561)) or
								((vState = 146) and (hState = 562)) or
								((vState = 146) and (hState = 565)) or
								((vState = 146) and (hState = 566)) or
								((vState = 146) and (hState = 567)) or
								((vState = 146) and (hState = 568)) or
								((vState = 146) and (hState = 572)) or
								((vState = 146) and (hState = 573)) or
								((vState = 146) and (hState = 574)) or
								((vState = 146) and (hState = 575)) or
								((vState = 146) and (hState = 576)) or
								((vState = 146) and (hState = 577)) or
								((vState = 146) and (hState = 578)) or
								((vState = 146) and (hState = 579)) or
								((vState = 146) and (hState = 580)) or
								((vState = 146) and (hState = 581)) or
								((vState = 146) and (hState = 582)) or
								((vState = 146) and (hState = 583)) or
								((vState = 146) and (hState = 584)) or
								((vState = 146) and (hState = 585)) or
								((vState = 146) and (hState = 586)) or
								((vState = 146) and (hState = 587)) or
								((vState = 146) and (hState = 588)) or
								((vState = 146) and (hState = 589)) or
								((vState = 146) and (hState = 590)) or
								((vState = 146) and (hState = 591)) or
								((vState = 146) and (hState = 592)) or
								((vState = 146) and (hState = 593)) or
								((vState = 146) and (hState = 594)) or
								((vState = 146) and (hState = 596)) or
								((vState = 146) and (hState = 597)) or
								((vState = 147) and (hState = 556)) or
								((vState = 147) and (hState = 557)) or
								((vState = 147) and (hState = 558)) or
								((vState = 147) and (hState = 561)) or
								((vState = 147) and (hState = 562)) or
								((vState = 147) and (hState = 565)) or
								((vState = 147) and (hState = 566)) or
								((vState = 147) and (hState = 567)) or
								((vState = 147) and (hState = 568)) or
								((vState = 147) and (hState = 572)) or
								((vState = 147) and (hState = 573)) or
								((vState = 147) and (hState = 574)) or
								((vState = 147) and (hState = 575)) or
								((vState = 147) and (hState = 579)) or
								((vState = 147) and (hState = 580)) or
								((vState = 147) and (hState = 581)) or
								((vState = 147) and (hState = 582)) or
								((vState = 147) and (hState = 583)) or
								((vState = 147) and (hState = 584)) or
								((vState = 147) and (hState = 585)) or
								((vState = 147) and (hState = 586)) or
								((vState = 147) and (hState = 587)) or
								((vState = 147) and (hState = 588)) or
								((vState = 147) and (hState = 589)) or
								((vState = 147) and (hState = 590)) or
								((vState = 147) and (hState = 591)) or
								((vState = 147) and (hState = 592)) or
								((vState = 147) and (hState = 593)) or
								((vState = 147) and (hState = 594)) or
								((vState = 147) and (hState = 595)) or
								((vState = 147) and (hState = 596)) or
								((vState = 147) and (hState = 597)) or
								((vState = 147) and (hState = 599)) or
								((vState = 148) and (hState = 557)) or
								((vState = 148) and (hState = 558)) or
								((vState = 148) and (hState = 562)) or
								((vState = 148) and (hState = 563)) or
								((vState = 148) and (hState = 565)) or
								((vState = 148) and (hState = 566)) or
								((vState = 148) and (hState = 567)) or
								((vState = 148) and (hState = 568)) or
								((vState = 148) and (hState = 569)) or
								((vState = 148) and (hState = 572)) or
								((vState = 148) and (hState = 573)) or
								((vState = 148) and (hState = 574)) or
								((vState = 148) and (hState = 577)) or
								((vState = 148) and (hState = 578)) or
								((vState = 148) and (hState = 579)) or
								((vState = 148) and (hState = 580)) or
								((vState = 148) and (hState = 581)) or
								((vState = 148) and (hState = 582)) or
								((vState = 148) and (hState = 583)) or
								((vState = 148) and (hState = 584)) or
								((vState = 148) and (hState = 585)) or
								((vState = 148) and (hState = 586)) or
								((vState = 148) and (hState = 587)) or
								((vState = 148) and (hState = 588)) or
								((vState = 148) and (hState = 589)) or
								((vState = 148) and (hState = 590)) or
								((vState = 148) and (hState = 591)) or
								((vState = 148) and (hState = 592)) or
								((vState = 148) and (hState = 593)) or
								((vState = 148) and (hState = 594)) or
								((vState = 148) and (hState = 595)) or
								((vState = 148) and (hState = 596)) or
								((vState = 148) and (hState = 599)) or
								((vState = 149) and (hState = 558)) or
								((vState = 149) and (hState = 559)) or
								((vState = 149) and (hState = 562)) or
								((vState = 149) and (hState = 563)) or
								((vState = 149) and (hState = 564)) or
								((vState = 149) and (hState = 566)) or
								((vState = 149) and (hState = 567)) or
								((vState = 149) and (hState = 568)) or
								((vState = 149) and (hState = 569)) or
								((vState = 149) and (hState = 570)) or
								((vState = 149) and (hState = 571)) or
								((vState = 149) and (hState = 572)) or
								((vState = 149) and (hState = 573)) or
								((vState = 149) and (hState = 574)) or
								((vState = 149) and (hState = 576)) or
								((vState = 149) and (hState = 577)) or
								((vState = 149) and (hState = 578)) or
								((vState = 149) and (hState = 582)) or
								((vState = 149) and (hState = 583)) or
								((vState = 149) and (hState = 584)) or
								((vState = 149) and (hState = 585)) or
								((vState = 149) and (hState = 586)) or
								((vState = 149) and (hState = 587)) or
								((vState = 149) and (hState = 588)) or
								((vState = 149) and (hState = 590)) or
								((vState = 149) and (hState = 591)) or
								((vState = 149) and (hState = 592)) or
								((vState = 149) and (hState = 593)) or
								((vState = 149) and (hState = 594)) or
								((vState = 149) and (hState = 595)) or
								((vState = 149) and (hState = 596)) or
								((vState = 149) and (hState = 599)) or
								((vState = 150) and (hState = 559)) or
								((vState = 150) and (hState = 560)) or
								((vState = 150) and (hState = 563)) or
								((vState = 150) and (hState = 564)) or
								((vState = 150) and (hState = 565)) or
								((vState = 150) and (hState = 566)) or
								((vState = 150) and (hState = 567)) or
								((vState = 150) and (hState = 569)) or
								((vState = 150) and (hState = 570)) or
								((vState = 150) and (hState = 571)) or
								((vState = 150) and (hState = 572)) or
								((vState = 150) and (hState = 573)) or
								((vState = 150) and (hState = 574)) or
								((vState = 150) and (hState = 575)) or
								((vState = 150) and (hState = 576)) or
								((vState = 150) and (hState = 577)) or
								((vState = 150) and (hState = 582)) or
								((vState = 150) and (hState = 583)) or
								((vState = 150) and (hState = 584)) or
								((vState = 150) and (hState = 585)) or
								((vState = 150) and (hState = 586)) or
								((vState = 150) and (hState = 587)) or
								((vState = 150) and (hState = 588)) or
								((vState = 150) and (hState = 589)) or
								((vState = 150) and (hState = 590)) or
								((vState = 150) and (hState = 591)) or
								((vState = 150) and (hState = 593)) or
								((vState = 150) and (hState = 594)) or
								((vState = 150) and (hState = 595)) or
								((vState = 150) and (hState = 596)) or
								((vState = 150) and (hState = 597)) or
								((vState = 150) and (hState = 599)) or
								((vState = 151) and (hState = 560)) or
								((vState = 151) and (hState = 561)) or
								((vState = 151) and (hState = 562)) or
								((vState = 151) and (hState = 563)) or
								((vState = 151) and (hState = 564)) or
								((vState = 151) and (hState = 565)) or
								((vState = 151) and (hState = 566)) or
								((vState = 151) and (hState = 567)) or
								((vState = 151) and (hState = 568)) or
								((vState = 151) and (hState = 569)) or
								((vState = 151) and (hState = 570)) or
								((vState = 151) and (hState = 571)) or
								((vState = 151) and (hState = 572)) or
								((vState = 151) and (hState = 573)) or
								((vState = 151) and (hState = 574)) or
								((vState = 151) and (hState = 575)) or
								((vState = 151) and (hState = 582)) or
								((vState = 151) and (hState = 583)) or
								((vState = 151) and (hState = 584)) or
								((vState = 151) and (hState = 585)) or
								((vState = 151) and (hState = 586)) or
								((vState = 151) and (hState = 587)) or
								((vState = 151) and (hState = 588)) or
								((vState = 151) and (hState = 589)) or
								((vState = 151) and (hState = 590)) or
								((vState = 151) and (hState = 592)) or
								((vState = 151) and (hState = 593)) or
								((vState = 151) and (hState = 594)) or
								((vState = 151) and (hState = 595)) or
								((vState = 151) and (hState = 596)) or
								((vState = 151) and (hState = 597)) or
								((vState = 151) and (hState = 598)) or
								((vState = 151) and (hState = 599)) or
								((vState = 152) and (hState = 562)) or
								((vState = 152) and (hState = 563)) or
								((vState = 152) and (hState = 564)) or
								((vState = 152) and (hState = 565)) or
								((vState = 152) and (hState = 566)) or
								((vState = 152) and (hState = 567)) or
								((vState = 152) and (hState = 568)) or
								((vState = 152) and (hState = 569)) or
								((vState = 152) and (hState = 570)) or
								((vState = 152) and (hState = 571)) or
								((vState = 152) and (hState = 572)) or
								((vState = 152) and (hState = 573)) or
								((vState = 152) and (hState = 574)) or
								((vState = 152) and (hState = 575)) or
								((vState = 152) and (hState = 581)) or
								((vState = 152) and (hState = 582)) or
								((vState = 152) and (hState = 583)) or
								((vState = 152) and (hState = 584)) or
								((vState = 152) and (hState = 585)) or
								((vState = 152) and (hState = 586)) or
								((vState = 152) and (hState = 587)) or
								((vState = 152) and (hState = 588)) or
								((vState = 152) and (hState = 589)) or
								((vState = 152) and (hState = 590)) or
								((vState = 152) and (hState = 591)) or
								((vState = 152) and (hState = 592)) or
								((vState = 152) and (hState = 593)) or
								((vState = 152) and (hState = 594)) or
								((vState = 152) and (hState = 597)) or
								((vState = 152) and (hState = 598)) or
								((vState = 152) and (hState = 599)) or
								((vState = 153) and (hState = 566)) or
								((vState = 153) and (hState = 567)) or
								((vState = 153) and (hState = 568)) or
								((vState = 153) and (hState = 569)) or
								((vState = 153) and (hState = 570)) or
								((vState = 153) and (hState = 571)) or
								((vState = 153) and (hState = 572)) or
								((vState = 153) and (hState = 573)) or
								((vState = 153) and (hState = 574)) or
								((vState = 153) and (hState = 575)) or
								((vState = 153) and (hState = 576)) or
								((vState = 153) and (hState = 577)) or
								((vState = 153) and (hState = 581)) or
								((vState = 153) and (hState = 582)) or
								((vState = 153) and (hState = 586)) or
								((vState = 153) and (hState = 587)) or
								((vState = 153) and (hState = 588)) or
								((vState = 153) and (hState = 589)) or
								((vState = 153) and (hState = 590)) or
								((vState = 153) and (hState = 591)) or
								((vState = 153) and (hState = 592)) or
								((vState = 153) and (hState = 593)) or
								((vState = 153) and (hState = 598)) or
								((vState = 154) and (hState = 567)) or
								((vState = 154) and (hState = 568)) or
								((vState = 154) and (hState = 573)) or
								((vState = 154) and (hState = 574)) or
								((vState = 154) and (hState = 575)) or
								((vState = 154) and (hState = 576)) or
								((vState = 154) and (hState = 577)) or
								((vState = 154) and (hState = 578)) or
								((vState = 154) and (hState = 579)) or
								((vState = 154) and (hState = 580)) or
								((vState = 154) and (hState = 581)) or
								((vState = 154) and (hState = 582)) or
								((vState = 154) and (hState = 587)) or
								((vState = 154) and (hState = 588)) or
								((vState = 154) and (hState = 589)) or
								((vState = 154) and (hState = 590)) or
								((vState = 154) and (hState = 591)) or
								((vState = 154) and (hState = 592)) or
								((vState = 154) and (hState = 593)) or
								((vState = 154) and (hState = 598)) or
								((vState = 154) and (hState = 599)) or
								((vState = 155) and (hState = 568)) or
								((vState = 155) and (hState = 569)) or
								((vState = 155) and (hState = 573)) or
								((vState = 155) and (hState = 574)) or
								((vState = 155) and (hState = 575)) or
								((vState = 155) and (hState = 576)) or
								((vState = 155) and (hState = 577)) or
								((vState = 155) and (hState = 578)) or
								((vState = 155) and (hState = 579)) or
								((vState = 155) and (hState = 580)) or
								((vState = 155) and (hState = 586)) or
								((vState = 155) and (hState = 587)) or
								((vState = 155) and (hState = 588)) or
								((vState = 155) and (hState = 589)) or
								((vState = 155) and (hState = 590)) or
								((vState = 155) and (hState = 591)) or
								((vState = 155) and (hState = 592)) or
								((vState = 155) and (hState = 598)) or
								((vState = 155) and (hState = 599)) or
								((vState = 156) and (hState = 568)) or
								((vState = 156) and (hState = 569)) or
								((vState = 156) and (hState = 570)) or
								((vState = 156) and (hState = 574)) or
								((vState = 156) and (hState = 575)) or
								((vState = 156) and (hState = 576)) or
								((vState = 156) and (hState = 577)) or
								((vState = 156) and (hState = 578)) or
								((vState = 156) and (hState = 579)) or
								((vState = 156) and (hState = 585)) or
								((vState = 156) and (hState = 586)) or
								((vState = 156) and (hState = 587)) or
								((vState = 156) and (hState = 589)) or
								((vState = 156) and (hState = 590)) or
								((vState = 156) and (hState = 591)) or
								((vState = 156) and (hState = 592)) or
								((vState = 156) and (hState = 598)) or
								((vState = 156) and (hState = 599)) or
								((vState = 157) and (hState = 569)) or
								((vState = 157) and (hState = 570)) or
								((vState = 157) and (hState = 571)) or
								((vState = 157) and (hState = 574)) or
								((vState = 157) and (hState = 575)) or
								((vState = 157) and (hState = 576)) or
								((vState = 157) and (hState = 577)) or
								((vState = 157) and (hState = 578)) or
								((vState = 157) and (hState = 579)) or
								((vState = 157) and (hState = 585)) or
								((vState = 157) and (hState = 586)) or
								((vState = 157) and (hState = 588)) or
								((vState = 157) and (hState = 589)) or
								((vState = 157) and (hState = 590)) or
								((vState = 157) and (hState = 591)) or
								((vState = 157) and (hState = 592)) or
								((vState = 157) and (hState = 593)) or
								((vState = 157) and (hState = 594)) or
								((vState = 157) and (hState = 598)) or
								((vState = 157) and (hState = 599)) or
								((vState = 158) and (hState = 570)) or
								((vState = 158) and (hState = 571)) or
								((vState = 158) and (hState = 574)) or
								((vState = 158) and (hState = 575)) or
								((vState = 158) and (hState = 576)) or
								((vState = 158) and (hState = 577)) or
								((vState = 158) and (hState = 578)) or
								((vState = 158) and (hState = 579)) or
								((vState = 158) and (hState = 580)) or
								((vState = 158) and (hState = 584)) or
								((vState = 158) and (hState = 585)) or
								((vState = 158) and (hState = 588)) or
								((vState = 158) and (hState = 589)) or
								((vState = 158) and (hState = 590)) or
								((vState = 158) and (hState = 591)) or
								((vState = 158) and (hState = 592)) or
								((vState = 158) and (hState = 593)) or
								((vState = 158) and (hState = 594)) or
								((vState = 158) and (hState = 595)) or
								((vState = 158) and (hState = 598)) or
								((vState = 158) and (hState = 599)) or
								((vState = 159) and (hState = 571)) or
								((vState = 159) and (hState = 572)) or
								((vState = 159) and (hState = 575)) or
								((vState = 159) and (hState = 576)) or
								((vState = 159) and (hState = 577)) or
								((vState = 159) and (hState = 579)) or
								((vState = 159) and (hState = 580)) or
								((vState = 159) and (hState = 581)) or
								((vState = 159) and (hState = 583)) or
								((vState = 159) and (hState = 584)) or
								((vState = 159) and (hState = 585)) or
								((vState = 159) and (hState = 587)) or
								((vState = 159) and (hState = 588)) or
								((vState = 159) and (hState = 591)) or
								((vState = 159) and (hState = 592)) or
								((vState = 159) and (hState = 593)) or
								((vState = 159) and (hState = 594)) or
								((vState = 159) and (hState = 595)) or
								((vState = 159) and (hState = 596)) or
								((vState = 159) and (hState = 598)) or
								((vState = 159) and (hState = 599)) or
								((vState = 160) and (hState = 572)) or
								((vState = 160) and (hState = 573)) or
								((vState = 160) and (hState = 576)) or
								((vState = 160) and (hState = 577)) or
								((vState = 160) and (hState = 580)) or
								((vState = 160) and (hState = 581)) or
								((vState = 160) and (hState = 582)) or
								((vState = 160) and (hState = 583)) or
								((vState = 160) and (hState = 584)) or
								((vState = 160) and (hState = 586)) or
								((vState = 160) and (hState = 587)) or
								((vState = 160) and (hState = 591)) or
								((vState = 160) and (hState = 592)) or
								((vState = 160) and (hState = 593)) or
								((vState = 160) and (hState = 595)) or
								((vState = 160) and (hState = 596)) or
								((vState = 160) and (hState = 597)) or
								((vState = 160) and (hState = 598)) or
								((vState = 160) and (hState = 599)) or
								((vState = 161) and (hState = 572)) or
								((vState = 161) and (hState = 573)) or
								((vState = 161) and (hState = 574)) or
								((vState = 161) and (hState = 577)) or
								((vState = 161) and (hState = 578)) or
								((vState = 161) and (hState = 581)) or
								((vState = 161) and (hState = 582)) or
								((vState = 161) and (hState = 583)) or
								((vState = 161) and (hState = 586)) or
								((vState = 161) and (hState = 587)) or
								((vState = 161) and (hState = 588)) or
								((vState = 161) and (hState = 591)) or
								((vState = 161) and (hState = 592)) or
								((vState = 161) and (hState = 593)) or
								((vState = 161) and (hState = 594)) or
								((vState = 161) and (hState = 596)) or
								((vState = 161) and (hState = 597)) or
								((vState = 161) and (hState = 598)) or
								((vState = 161) and (hState = 599)) or
								((vState = 162) and (hState = 573)) or
								((vState = 162) and (hState = 574)) or
								((vState = 162) and (hState = 575)) or
								((vState = 162) and (hState = 578)) or
								((vState = 162) and (hState = 579)) or
								((vState = 162) and (hState = 581)) or
								((vState = 162) and (hState = 582)) or
								((vState = 162) and (hState = 583)) or
								((vState = 162) and (hState = 584)) or
								((vState = 162) and (hState = 587)) or
								((vState = 162) and (hState = 588)) or
								((vState = 162) and (hState = 591)) or
								((vState = 162) and (hState = 592)) or
								((vState = 162) and (hState = 593)) or
								((vState = 162) and (hState = 594)) or
								((vState = 162) and (hState = 597)) or
								((vState = 162) and (hState = 598)) or
								((vState = 162) and (hState = 599)) or
								((vState = 163) and (hState = 574)) or
								((vState = 163) and (hState = 575)) or
								((vState = 163) and (hState = 578)) or
								((vState = 163) and (hState = 579)) or
								((vState = 163) and (hState = 580)) or
								((vState = 163) and (hState = 581)) or
								((vState = 163) and (hState = 582)) or
								((vState = 163) and (hState = 583)) or
								((vState = 163) and (hState = 584)) or
								((vState = 163) and (hState = 585)) or
								((vState = 163) and (hState = 588)) or
								((vState = 163) and (hState = 589)) or
								((vState = 163) and (hState = 590)) or
								((vState = 163) and (hState = 591)) or
								((vState = 163) and (hState = 592)) or
								((vState = 163) and (hState = 593)) or
								((vState = 163) and (hState = 594)) or
								((vState = 163) and (hState = 595)) or
								((vState = 163) and (hState = 596)) or
								((vState = 163) and (hState = 597)) or
								((vState = 163) and (hState = 598)) or
								((vState = 163) and (hState = 599)) or
								((vState = 164) and (hState = 575)) or
								((vState = 164) and (hState = 576)) or
								((vState = 164) and (hState = 579)) or
								((vState = 164) and (hState = 580)) or
								((vState = 164) and (hState = 581)) or
								((vState = 164) and (hState = 584)) or
								((vState = 164) and (hState = 585)) or
								((vState = 164) and (hState = 586)) or
								((vState = 164) and (hState = 588)) or
								((vState = 164) and (hState = 589)) or
								((vState = 164) and (hState = 590)) or
								((vState = 164) and (hState = 591)) or
								((vState = 164) and (hState = 592)) or
								((vState = 164) and (hState = 593)) or
								((vState = 164) and (hState = 594)) or
								((vState = 164) and (hState = 595)) or
								((vState = 164) and (hState = 596)) or
								((vState = 164) and (hState = 597)) or
								((vState = 164) and (hState = 599)) or
								((vState = 165) and (hState = 576)) or
								((vState = 165) and (hState = 577)) or
								((vState = 165) and (hState = 579)) or
								((vState = 165) and (hState = 580)) or
								((vState = 165) and (hState = 581)) or
								((vState = 165) and (hState = 585)) or
								((vState = 165) and (hState = 586)) or
								((vState = 165) and (hState = 587)) or
								((vState = 165) and (hState = 589)) or
								((vState = 165) and (hState = 590)) or
								((vState = 165) and (hState = 591)) or
								((vState = 165) and (hState = 592)) or
								((vState = 165) and (hState = 593)) or
								((vState = 165) and (hState = 594)) or
								((vState = 165) and (hState = 595)) or
								((vState = 165) and (hState = 596)) or
								((vState = 165) and (hState = 597)) or
								((vState = 165) and (hState = 599)) or
								((vState = 166) and (hState = 577)) or
								((vState = 166) and (hState = 578)) or
								((vState = 166) and (hState = 579)) or
								((vState = 166) and (hState = 580)) or
								((vState = 166) and (hState = 581)) or
								((vState = 166) and (hState = 586)) or
								((vState = 166) and (hState = 587)) or
								((vState = 166) and (hState = 589)) or
								((vState = 166) and (hState = 590)) or
								((vState = 166) and (hState = 591)) or
								((vState = 166) and (hState = 592)) or
								((vState = 166) and (hState = 593)) or
								((vState = 166) and (hState = 594)) or
								((vState = 166) and (hState = 595)) or
								((vState = 166) and (hState = 596)) or
								((vState = 166) and (hState = 597)) or
								((vState = 166) and (hState = 598)) or
								((vState = 166) and (hState = 599)) or
								((vState = 167) and (hState = 577)) or
								((vState = 167) and (hState = 578)) or
								((vState = 167) and (hState = 579)) or
								((vState = 167) and (hState = 581)) or
								((vState = 167) and (hState = 582)) or
								((vState = 167) and (hState = 586)) or
								((vState = 167) and (hState = 587)) or
								((vState = 167) and (hState = 590)) or
								((vState = 167) and (hState = 591)) or
								((vState = 167) and (hState = 592)) or
								((vState = 167) and (hState = 593)) or
								((vState = 167) and (hState = 594)) or
								((vState = 167) and (hState = 595)) or
								((vState = 167) and (hState = 596)) or
								((vState = 167) and (hState = 597)) or
								((vState = 167) and (hState = 598)) or
								((vState = 167) and (hState = 599)) or
								((vState = 168) and (hState = 577)) or
								((vState = 168) and (hState = 578)) or
								((vState = 168) and (hState = 579)) or
								((vState = 168) and (hState = 581)) or
								((vState = 168) and (hState = 582)) or
								((vState = 168) and (hState = 583)) or
								((vState = 168) and (hState = 586)) or
								((vState = 168) and (hState = 587)) or
								((vState = 168) and (hState = 589)) or
								((vState = 168) and (hState = 590)) or
								((vState = 168) and (hState = 591)) or
								((vState = 168) and (hState = 592)) or
								((vState = 168) and (hState = 593)) or
								((vState = 168) and (hState = 594)) or
								((vState = 168) and (hState = 595)) or
								((vState = 168) and (hState = 596)) or
								((vState = 168) and (hState = 597)) or
								((vState = 168) and (hState = 598)) or
								((vState = 168) and (hState = 599)) or
								((vState = 169) and (hState = 576)) or
								((vState = 169) and (hState = 577)) or
								((vState = 169) and (hState = 578)) or
								((vState = 169) and (hState = 582)) or
								((vState = 169) and (hState = 583)) or
								((vState = 169) and (hState = 586)) or
								((vState = 169) and (hState = 587)) or
								((vState = 169) and (hState = 588)) or
								((vState = 169) and (hState = 589)) or
								((vState = 169) and (hState = 590)) or
								((vState = 169) and (hState = 591)) or
								((vState = 169) and (hState = 592)) or
								((vState = 169) and (hState = 593)) or
								((vState = 169) and (hState = 594)) or
								((vState = 169) and (hState = 595)) or
								((vState = 169) and (hState = 596)) or
								((vState = 169) and (hState = 598)) or
								((vState = 169) and (hState = 599)) or
								((vState = 170) and (hState = 575)) or
								((vState = 170) and (hState = 576)) or
								((vState = 170) and (hState = 577)) or
								((vState = 170) and (hState = 578)) or
								((vState = 170) and (hState = 583)) or
								((vState = 170) and (hState = 584)) or
								((vState = 170) and (hState = 585)) or
								((vState = 170) and (hState = 586)) or
								((vState = 170) and (hState = 587)) or
								((vState = 170) and (hState = 588)) or
								((vState = 170) and (hState = 589)) or
								((vState = 170) and (hState = 590)) or
								((vState = 170) and (hState = 591)) or
								((vState = 170) and (hState = 592)) or
								((vState = 170) and (hState = 593)) or
								((vState = 170) and (hState = 594)) or
								((vState = 170) and (hState = 595)) or
								((vState = 170) and (hState = 599)) or
								((vState = 171) and (hState = 574)) or
								((vState = 171) and (hState = 575)) or
								((vState = 171) and (hState = 576)) or
								((vState = 171) and (hState = 577)) or
								((vState = 171) and (hState = 582)) or
								((vState = 171) and (hState = 583)) or
								((vState = 171) and (hState = 584)) or
								((vState = 171) and (hState = 585)) or
								((vState = 171) and (hState = 586)) or
								((vState = 171) and (hState = 587)) or
								((vState = 171) and (hState = 588)) or
								((vState = 171) and (hState = 589)) or
								((vState = 171) and (hState = 590)) or
								((vState = 171) and (hState = 591)) or
								((vState = 171) and (hState = 592)) or
								((vState = 171) and (hState = 593)) or
								((vState = 171) and (hState = 594)) or
								((vState = 171) and (hState = 595)) or
								((vState = 172) and (hState = 574)) or
								((vState = 172) and (hState = 575)) or
								((vState = 172) and (hState = 576)) or
								((vState = 172) and (hState = 579)) or
								((vState = 172) and (hState = 580)) or
								((vState = 172) and (hState = 581)) or
								((vState = 172) and (hState = 582)) or
								((vState = 172) and (hState = 583)) or
								((vState = 172) and (hState = 584)) or
								((vState = 172) and (hState = 585)) or
								((vState = 172) and (hState = 586)) or
								((vState = 172) and (hState = 587)) or
								((vState = 172) and (hState = 588)) or
								((vState = 172) and (hState = 589)) or
								((vState = 172) and (hState = 590)) or
								((vState = 172) and (hState = 591)) or
								((vState = 172) and (hState = 592)) or
								((vState = 172) and (hState = 593)) or
								((vState = 172) and (hState = 594)) or
								((vState = 172) and (hState = 595)) or
								((vState = 172) and (hState = 596)) or
								((vState = 173) and (hState = 573)) or
								((vState = 173) and (hState = 574)) or
								((vState = 173) and (hState = 575)) or
								((vState = 173) and (hState = 576)) or
								((vState = 173) and (hState = 578)) or
								((vState = 173) and (hState = 579)) or
								((vState = 173) and (hState = 580)) or
								((vState = 173) and (hState = 581)) or
								((vState = 173) and (hState = 585)) or
								((vState = 173) and (hState = 586)) or
								((vState = 173) and (hState = 587)) or
								((vState = 173) and (hState = 588)) or
								((vState = 173) and (hState = 589)) or
								((vState = 173) and (hState = 590)) or
								((vState = 173) and (hState = 591)) or
								((vState = 173) and (hState = 592)) or
								((vState = 173) and (hState = 593)) or
								((vState = 173) and (hState = 594)) or
								((vState = 173) and (hState = 595)) or
								((vState = 173) and (hState = 596)) or
								((vState = 174) and (hState = 573)) or
								((vState = 174) and (hState = 574)) or
								((vState = 174) and (hState = 575)) or
								((vState = 174) and (hState = 579)) or
								((vState = 174) and (hState = 580)) or
								((vState = 174) and (hState = 585)) or
								((vState = 174) and (hState = 586)) or
								((vState = 174) and (hState = 587)) or
								((vState = 174) and (hState = 591)) or
								((vState = 174) and (hState = 592)) or
								((vState = 174) and (hState = 593)) or
								((vState = 174) and (hState = 594)) or
								((vState = 174) and (hState = 595)) or
								((vState = 174) and (hState = 596)) or
								((vState = 175) and (hState = 573)) or
								((vState = 175) and (hState = 574)) or
								((vState = 175) and (hState = 575)) or
								((vState = 175) and (hState = 576)) or
								((vState = 175) and (hState = 580)) or
								((vState = 175) and (hState = 581)) or
								((vState = 175) and (hState = 582)) or
								((vState = 175) and (hState = 584)) or
								((vState = 175) and (hState = 585)) or
								((vState = 175) and (hState = 586)) or
								((vState = 175) and (hState = 587)) or
								((vState = 175) and (hState = 592)) or
								((vState = 175) and (hState = 593)) or
								((vState = 175) and (hState = 594)) or
								((vState = 175) and (hState = 595)) or
								((vState = 175) and (hState = 596)) or
								((vState = 175) and (hState = 597)) or
								((vState = 175) and (hState = 598)) or
								((vState = 175) and (hState = 599)) or
								((vState = 176) and (hState = 575)) or
								((vState = 176) and (hState = 576)) or
								((vState = 176) and (hState = 577)) or
								((vState = 176) and (hState = 581)) or
								((vState = 176) and (hState = 582)) or
								((vState = 176) and (hState = 583)) or
								((vState = 176) and (hState = 584)) or
								((vState = 176) and (hState = 585)) or
								((vState = 176) and (hState = 586)) or
								((vState = 176) and (hState = 592)) or
								((vState = 176) and (hState = 593)) or
								((vState = 176) and (hState = 594)) or
								((vState = 176) and (hState = 595)) or
								((vState = 176) and (hState = 596)) or
								((vState = 176) and (hState = 597)) or
								((vState = 176) and (hState = 598)) or
								((vState = 176) and (hState = 599)) or
								((vState = 177) and (hState = 577)) or
								((vState = 177) and (hState = 578)) or
								((vState = 177) and (hState = 579)) or
								((vState = 177) and (hState = 582)) or
								((vState = 177) and (hState = 583)) or
								((vState = 177) and (hState = 584)) or
								((vState = 177) and (hState = 585)) or
								((vState = 177) and (hState = 586)) or
								((vState = 177) and (hState = 592)) or
								((vState = 177) and (hState = 593)) or
								((vState = 177) and (hState = 594)) or
								((vState = 177) and (hState = 595)) or
								((vState = 177) and (hState = 596)) or
								((vState = 177) and (hState = 597)) or
								((vState = 177) and (hState = 599)) or
								((vState = 178) and (hState = 578)) or
								((vState = 178) and (hState = 579)) or
								((vState = 178) and (hState = 580)) or
								((vState = 178) and (hState = 581)) or
								((vState = 178) and (hState = 584)) or
								((vState = 178) and (hState = 585)) or
								((vState = 178) and (hState = 590)) or
								((vState = 178) and (hState = 591)) or
								((vState = 178) and (hState = 592)) or
								((vState = 178) and (hState = 593)) or
								((vState = 178) and (hState = 594)) or
								((vState = 178) and (hState = 595)) or
								((vState = 178) and (hState = 596)) or
								((vState = 178) and (hState = 597)) or
								((vState = 179) and (hState = 580)) or
								((vState = 179) and (hState = 581)) or
								((vState = 179) and (hState = 582)) or
								((vState = 179) and (hState = 584)) or
								((vState = 179) and (hState = 585)) or
								((vState = 179) and (hState = 586)) or
								((vState = 179) and (hState = 587)) or
								((vState = 179) and (hState = 589)) or
								((vState = 179) and (hState = 590)) or
								((vState = 179) and (hState = 591)) or
								((vState = 179) and (hState = 592)) or
								((vState = 179) and (hState = 593)) or
								((vState = 179) and (hState = 594)) or
								((vState = 179) and (hState = 596)) or
								((vState = 179) and (hState = 597)) or
								((vState = 179) and (hState = 598)) or
								((vState = 180) and (hState = 581)) or
								((vState = 180) and (hState = 582)) or
								((vState = 180) and (hState = 583)) or
								((vState = 180) and (hState = 585)) or
								((vState = 180) and (hState = 586)) or
								((vState = 180) and (hState = 587)) or
								((vState = 180) and (hState = 588)) or
								((vState = 180) and (hState = 589)) or
								((vState = 180) and (hState = 590)) or
								((vState = 180) and (hState = 591)) or
								((vState = 180) and (hState = 592)) or
								((vState = 180) and (hState = 593)) or
								((vState = 180) and (hState = 594)) or
								((vState = 180) and (hState = 596)) or
								((vState = 180) and (hState = 597)) or
								((vState = 180) and (hState = 598)) or
								((vState = 181) and (hState = 583)) or
								((vState = 181) and (hState = 584)) or
								((vState = 181) and (hState = 585)) or
								((vState = 181) and (hState = 586)) or
								((vState = 181) and (hState = 587)) or
								((vState = 181) and (hState = 588)) or
								((vState = 181) and (hState = 589)) or
								((vState = 181) and (hState = 590)) or
								((vState = 181) and (hState = 591)) or
								((vState = 181) and (hState = 592)) or
								((vState = 181) and (hState = 593)) or
								((vState = 181) and (hState = 594)) or
								((vState = 181) and (hState = 597)) or
								((vState = 181) and (hState = 598)) or
								((vState = 182) and (hState = 584)) or
								((vState = 182) and (hState = 585)) or
								((vState = 182) and (hState = 586)) or
								((vState = 182) and (hState = 587)) or
								((vState = 182) and (hState = 588)) or
								((vState = 182) and (hState = 589)) or
								((vState = 182) and (hState = 590)) or
								((vState = 182) and (hState = 592)) or
								((vState = 182) and (hState = 593)) or
								((vState = 182) and (hState = 594)) or
								((vState = 183) and (hState = 586)) or
								((vState = 183) and (hState = 587)) or
								((vState = 183) and (hState = 588)) or
								((vState = 183) and (hState = 589)) or
								((vState = 183) and (hState = 590)) or
								((vState = 183) and (hState = 591)) or
								((vState = 183) and (hState = 593)) or
								((vState = 183) and (hState = 594)) or
								((vState = 183) and (hState = 595)) or
								((vState = 183) and (hState = 596)) or
								((vState = 184) and (hState = 587)) or
								((vState = 184) and (hState = 588)) or
								((vState = 184) and (hState = 589)) or
								((vState = 184) and (hState = 590)) or
								((vState = 184) and (hState = 591)) or
								((vState = 184) and (hState = 592)) or
								((vState = 184) and (hState = 593)) or
								((vState = 184) and (hState = 594)) or
								((vState = 184) and (hState = 595)) or
								((vState = 184) and (hState = 596)) or
								((vState = 184) and (hState = 597)) or
								((vState = 185) and (hState = 589)) or
								((vState = 185) and (hState = 590)) or
								((vState = 185) and (hState = 591)) or
								((vState = 185) and (hState = 592)) or
								((vState = 185) and (hState = 593)) or
								((vState = 185) and (hState = 594)) or
								((vState = 185) and (hState = 596)) or
								((vState = 185) and (hState = 597)) or
								((vState = 185) and (hState = 598)) or
								((vState = 186) and (hState = 590)) or
								((vState = 186) and (hState = 591)) or
								((vState = 186) and (hState = 593)) or
								((vState = 186) and (hState = 594)) or
								((vState = 186) and (hState = 595)) or
								((vState = 186) and (hState = 598)) or
								((vState = 186) and (hState = 599)) or
								((vState = 187) and (hState = 591)) or
								((vState = 187) and (hState = 592)) or
								((vState = 187) and (hState = 594)) or
								((vState = 187) and (hState = 599)) or
								((vState = 188) and (hState = 591)) or
								((vState = 188) and (hState = 592)) or
								((vState = 188) and (hState = 593)) or
								((vState = 189) and (hState = 592)) or
								((vState = 189) and (hState = 593)) or
								((vState = 189) and (hState = 594)) or
								((vState = 190) and (hState = 593)) or
								((vState = 190) and (hState = 594)) or
								((vState = 190) and (hState = 595)) or
								((vState = 191) and (hState = 594)) or
								((vState = 191) and (hState = 595)) else (others => '0');
end architecture me;

library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity picture is
	port (
		vState : in std_logic_vector(15 downto 0);
		hState : in std_logic_vector(15 downto 0);
		r : out std_logic;
		g : out std_logic;
		b : out std_logic
	);
end entity picture;

architecture first of picture is
	
begin
	r <= '1' when vState < 100 else '0';
	g <= '1' when hState > 300 else '0';
	b <= '1' when vState * vState < 300*400 else '0';
	
end architecture first;

architecture me of picture is
	signal rgb : std_logic_vector(2 downto 0);
	
begin
	r <= rgb(0);
	g <= rgb(1);
	b <= rgb(2);
	
	rgb <= (others => '1') when ((vState = 176) and (hState = 578)) or
								((vState = 176) and (hState = 579)) or
								((vState = 176) and (hState = 587)) or
								((vState = 176) and (hState = 588)) or
								((vState = 176) and (hState = 589)) or
								((vState = 176) and (hState = 590)) or
								((vState = 176) and (hState = 591)) or
								((vState = 176) and (hState = 592)) or
								((vState = 176) and (hState = 593)) or
								((vState = 177) and (hState = 578)) or
								((vState = 177) and (hState = 579)) or
								((vState = 177) and (hState = 587)) or
								((vState = 177) and (hState = 588)) or
								((vState = 177) and (hState = 589)) or
								((vState = 177) and (hState = 590)) or
								((vState = 177) and (hState = 591)) or
								((vState = 177) and (hState = 592)) or
								((vState = 177) and (hState = 593)) or
								((vState = 178) and (hState = 595)) or
								((vState = 178) and (hState = 596)) or
								((vState = 178) and (hState = 597)) or
								((vState = 178) and (hState = 598)) or
								((vState = 178) and (hState = 599)) or
								((vState = 182) and (hState = 584)) or
								((vState = 183) and (hState = 585)) or
								((vState = 184) and (hState = 588)) or
								((vState = 184) and (hState = 595)) or
								((vState = 187) and (hState = 590)) or
								((vState = 187) and (hState = 591)) or
								((vState = 188) and (hState = 590)) or
								((vState = 188) and (hState = 591)) or
								((vState = 189) and (hState = 588)) or
								((vState = 190) and (hState = 595)) or
								((vState = 192) and (hState = 584)) or
								((vState = 193) and (hState = 583)) or
								((vState = 193) and (hState = 584)) or
								((vState = 194) and (hState = 581)) or
								((vState = 194) and (hState = 582)) or
								((vState = 194) and (hState = 583)) or
								((vState = 194) and (hState = 595)) or
								((vState = 195) and (hState = 579)) or
								((vState = 195) and (hState = 580)) or
								((vState = 195) and (hState = 581)) or
								((vState = 196) and (hState = 579)) or
								((vState = 196) and (hState = 580)) or
								((vState = 197) and (hState = 578)) or
								((vState = 197) and (hState = 579)) or
								((vState = 198) and (hState = 576)) or
								((vState = 198) and (hState = 577)) or
								((vState = 198) and (hState = 578)) or
								((vState = 198) and (hState = 579)) or
								((vState = 198) and (hState = 593)) or
								((vState = 199) and (hState = 574)) or
								((vState = 199) and (hState = 575)) or
								((vState = 199) and (hState = 576)) or
								((vState = 199) and (hState = 577)) or
								((vState = 199) and (hState = 578)) or
								((vState = 200) and (hState = 572)) or
								((vState = 200) and (hState = 576)) or
								((vState = 200) and (hState = 577)) or
								((vState = 200) and (hState = 590)) or
								((vState = 205) and (hState = 547)) or
								((vState = 206) and (hState = 548)) or
								((vState = 206) and (hState = 559)) or
								((vState = 209) and (hState = 551)) or
								((vState = 209) and (hState = 561)) or
								((vState = 209) and (hState = 567)) or
								((vState = 209) and (hState = 583)) or
								((vState = 210) and (hState = 551)) or
								((vState = 210) and (hState = 552)) or
								((vState = 210) and (hState = 553)) or
								((vState = 210) and (hState = 562)) or
								((vState = 211) and (hState = 551)) or
								((vState = 211) and (hState = 552)) or
								((vState = 211) and (hState = 553)) or
								((vState = 211) and (hState = 563)) or
								((vState = 211) and (hState = 564)) or
								((vState = 212) and (hState = 563)) or
								((vState = 212) and (hState = 564)) or
								((vState = 213) and (hState = 563)) or
								((vState = 213) and (hState = 564)) or
								((vState = 214) and (hState = 548)) or
								((vState = 214) and (hState = 556)) or
								((vState = 214) and (hState = 562)) or
								((vState = 214) and (hState = 563)) or
								((vState = 214) and (hState = 564)) or
								((vState = 214) and (hState = 579)) or
								((vState = 214) and (hState = 594)) or
								((vState = 214) and (hState = 595)) or
								((vState = 214) and (hState = 596)) or
								((vState = 215) and (hState = 544)) or
								((vState = 215) and (hState = 545)) or
								((vState = 215) and (hState = 546)) or
								((vState = 215) and (hState = 547)) or
								((vState = 215) and (hState = 557)) or
								((vState = 215) and (hState = 578)) or
								((vState = 215) and (hState = 589)) or
								((vState = 215) and (hState = 590)) or
								((vState = 215) and (hState = 591)) or
								((vState = 215) and (hState = 592)) or
								((vState = 215) and (hState = 593)) or
								((vState = 215) and (hState = 594)) or
								((vState = 216) and (hState = 542)) or
								((vState = 216) and (hState = 543)) or
								((vState = 216) and (hState = 544)) or
								((vState = 216) and (hState = 545)) or
								((vState = 216) and (hState = 546)) or
								((vState = 216) and (hState = 547)) or
								((vState = 216) and (hState = 558)) or
								((vState = 216) and (hState = 559)) or
								((vState = 216) and (hState = 560)) or
								((vState = 216) and (hState = 567)) or
								((vState = 216) and (hState = 584)) or
								((vState = 216) and (hState = 585)) or
								((vState = 216) and (hState = 586)) or
								((vState = 216) and (hState = 590)) or
								((vState = 216) and (hState = 591)) or
								((vState = 217) and (hState = 542)) or
								((vState = 217) and (hState = 543)) or
								((vState = 217) and (hState = 558)) or
								((vState = 217) and (hState = 559)) or
								((vState = 217) and (hState = 560)) or
								((vState = 217) and (hState = 590)) or
								((vState = 218) and (hState = 541)) or
								((vState = 218) and (hState = 558)) or
								((vState = 218) and (hState = 559)) or
								((vState = 218) and (hState = 560)) or
								((vState = 218) and (hState = 561)) or
								((vState = 218) and (hState = 577)) or
								((vState = 219) and (hState = 539)) or
								((vState = 219) and (hState = 540)) or
								((vState = 219) and (hState = 541)) or
								((vState = 219) and (hState = 552)) or
								((vState = 219) and (hState = 558)) or
								((vState = 219) and (hState = 559)) or
								((vState = 219) and (hState = 560)) or
								((vState = 219) and (hState = 561)) or
								((vState = 219) and (hState = 562)) or
								((vState = 219) and (hState = 568)) or
								((vState = 219) and (hState = 576)) or
								((vState = 219) and (hState = 577)) or
								((vState = 219) and (hState = 578)) or
								((vState = 219) and (hState = 588)) or
								((vState = 220) and (hState = 537)) or
								((vState = 220) and (hState = 538)) or
								((vState = 220) and (hState = 539)) or
								((vState = 220) and (hState = 540)) or
								((vState = 220) and (hState = 558)) or
								((vState = 220) and (hState = 559)) or
								((vState = 220) and (hState = 560)) or
								((vState = 220) and (hState = 561)) or
								((vState = 220) and (hState = 562)) or
								((vState = 220) and (hState = 563)) or
								((vState = 220) and (hState = 569)) or
								((vState = 220) and (hState = 570)) or
								((vState = 220) and (hState = 571)) or
								((vState = 220) and (hState = 572)) or
								((vState = 220) and (hState = 573)) or
								((vState = 220) and (hState = 574)) or
								((vState = 220) and (hState = 585)) or
								((vState = 221) and (hState = 536)) or
								((vState = 221) and (hState = 537)) or
								((vState = 221) and (hState = 557)) or
								((vState = 221) and (hState = 558)) or
								((vState = 221) and (hState = 559)) or
								((vState = 221) and (hState = 560)) or
								((vState = 221) and (hState = 561)) or
								((vState = 221) and (hState = 562)) or
								((vState = 221) and (hState = 563)) or
								((vState = 221) and (hState = 564)) or
								((vState = 221) and (hState = 569)) or
								((vState = 221) and (hState = 570)) or
								((vState = 221) and (hState = 571)) or
								((vState = 221) and (hState = 572)) or
								((vState = 221) and (hState = 573)) or
								((vState = 221) and (hState = 585)) or
								((vState = 222) and (hState = 536)) or
								((vState = 222) and (hState = 560)) or
								((vState = 222) and (hState = 561)) or
								((vState = 222) and (hState = 562)) or
								((vState = 222) and (hState = 563)) or
								((vState = 222) and (hState = 564)) or
								((vState = 222) and (hState = 565)) or
								((vState = 222) and (hState = 569)) or
								((vState = 222) and (hState = 570)) or
								((vState = 222) and (hState = 571)) or
								((vState = 222) and (hState = 572)) or
								((vState = 222) and (hState = 585)) or
								((vState = 223) and (hState = 535)) or
								((vState = 223) and (hState = 561)) or
								((vState = 223) and (hState = 562)) or
								((vState = 223) and (hState = 563)) or
								((vState = 223) and (hState = 564)) or
								((vState = 223) and (hState = 565)) or
								((vState = 223) and (hState = 566)) or
								((vState = 223) and (hState = 569)) or
								((vState = 223) and (hState = 570)) or
								((vState = 223) and (hState = 571)) or
								((vState = 223) and (hState = 572)) or
								((vState = 223) and (hState = 585)) or
								((vState = 224) and (hState = 563)) or
								((vState = 224) and (hState = 564)) or
								((vState = 224) and (hState = 565)) or
								((vState = 224) and (hState = 566)) or
								((vState = 224) and (hState = 567)) or
								((vState = 224) and (hState = 568)) or
								((vState = 224) and (hState = 569)) or
								((vState = 224) and (hState = 570)) or
								((vState = 224) and (hState = 571)) or
								((vState = 224) and (hState = 572)) or
								((vState = 225) and (hState = 532)) or
								((vState = 225) and (hState = 563)) or
								((vState = 225) and (hState = 564)) or
								((vState = 225) and (hState = 565)) or
								((vState = 225) and (hState = 566)) or
								((vState = 225) and (hState = 567)) or
								((vState = 225) and (hState = 568)) or
								((vState = 225) and (hState = 569)) or
								((vState = 225) and (hState = 570)) or
								((vState = 225) and (hState = 571)) or
								((vState = 225) and (hState = 572)) or
								((vState = 225) and (hState = 573)) or
								((vState = 226) and (hState = 530)) or
								((vState = 226) and (hState = 531)) or
								((vState = 226) and (hState = 566)) or
								((vState = 226) and (hState = 567)) or
								((vState = 226) and (hState = 568)) or
								((vState = 226) and (hState = 569)) or
								((vState = 226) and (hState = 570)) or
								((vState = 226) and (hState = 574)) or
								((vState = 227) and (hState = 529)) or
								((vState = 227) and (hState = 530)) or
								((vState = 227) and (hState = 568)) or
								((vState = 227) and (hState = 569)) or
								((vState = 227) and (hState = 570)) or
								((vState = 227) and (hState = 574)) or
								((vState = 228) and (hState = 568)) or
								((vState = 228) and (hState = 569)) or
								((vState = 228) and (hState = 570)) or
								((vState = 228) and (hState = 571)) or
								((vState = 228) and (hState = 574)) or
								((vState = 229) and (hState = 568)) or
								((vState = 229) and (hState = 569)) or
								((vState = 229) and (hState = 570)) or
								((vState = 229) and (hState = 571)) or
								((vState = 229) and (hState = 572)) or
								((vState = 229) and (hState = 573)) or
								((vState = 229) and (hState = 574)) or
								((vState = 229) and (hState = 575)) or
								((vState = 230) and (hState = 567)) or
								((vState = 230) and (hState = 568)) or
								((vState = 230) and (hState = 569)) or
								((vState = 230) and (hState = 570)) or
								((vState = 230) and (hState = 571)) or
								((vState = 230) and (hState = 572)) or
								((vState = 230) and (hState = 573)) or
								((vState = 230) and (hState = 574)) or
								((vState = 230) and (hState = 575)) or
								((vState = 230) and (hState = 576)) or
								((vState = 230) and (hState = 577)) or
								((vState = 231) and (hState = 566)) or
								((vState = 231) and (hState = 567)) or
								((vState = 231) and (hState = 568)) or
								((vState = 231) and (hState = 572)) or
								((vState = 231) and (hState = 573)) or
								((vState = 231) and (hState = 574)) or
								((vState = 231) and (hState = 575)) or
								((vState = 231) and (hState = 576)) or
								((vState = 231) and (hState = 577)) or
								((vState = 231) and (hState = 588)) or
								((vState = 232) and (hState = 565)) or
								((vState = 232) and (hState = 566)) or
								((vState = 232) and (hState = 567)) or
								((vState = 232) and (hState = 573)) or
								((vState = 232) and (hState = 574)) or
								((vState = 232) and (hState = 575)) or
								((vState = 232) and (hState = 576)) or
								((vState = 232) and (hState = 577)) or
								((vState = 232) and (hState = 578)) or
								((vState = 232) and (hState = 588)) or
								((vState = 233) and (hState = 567)) or
								((vState = 233) and (hState = 574)) or
								((vState = 233) and (hState = 575)) or
								((vState = 233) and (hState = 576)) or
								((vState = 233) and (hState = 577)) or
								((vState = 233) and (hState = 578)) or
								((vState = 233) and (hState = 588)) or
								((vState = 234) and (hState = 567)) or
								((vState = 234) and (hState = 574)) or
								((vState = 234) and (hState = 575)) or
								((vState = 234) and (hState = 576)) or
								((vState = 234) and (hState = 577)) or
								((vState = 234) and (hState = 578)) or
								((vState = 234) and (hState = 579)) or
								((vState = 234) and (hState = 580)) or
								((vState = 234) and (hState = 584)) or
								((vState = 234) and (hState = 585)) or
								((vState = 234) and (hState = 586)) or
								((vState = 234) and (hState = 587)) or
								((vState = 234) and (hState = 588)) or
								((vState = 234) and (hState = 589)) or
								((vState = 234) and (hState = 590)) or
								((vState = 235) and (hState = 567)) or
								((vState = 235) and (hState = 574)) or
								((vState = 235) and (hState = 575)) or
								((vState = 235) and (hState = 576)) or
								((vState = 235) and (hState = 577)) or
								((vState = 235) and (hState = 578)) or
								((vState = 235) and (hState = 579)) or
								((vState = 235) and (hState = 580)) or
								((vState = 235) and (hState = 581)) or
								((vState = 235) and (hState = 582)) or
								((vState = 235) and (hState = 583)) or
								((vState = 235) and (hState = 584)) or
								((vState = 235) and (hState = 585)) or
								((vState = 235) and (hState = 586)) or
								((vState = 235) and (hState = 587)) or
								((vState = 235) and (hState = 588)) or
								((vState = 235) and (hState = 589)) or
								((vState = 235) and (hState = 590)) or
								((vState = 236) and (hState = 562)) or
								((vState = 236) and (hState = 567)) or
								((vState = 236) and (hState = 568)) or
								((vState = 236) and (hState = 569)) or
								((vState = 236) and (hState = 570)) or
								((vState = 236) and (hState = 571)) or
								((vState = 236) and (hState = 572)) or
								((vState = 236) and (hState = 573)) or
								((vState = 236) and (hState = 574)) or
								((vState = 236) and (hState = 575)) or
								((vState = 236) and (hState = 576)) or
								((vState = 236) and (hState = 577)) or
								((vState = 236) and (hState = 578)) or
								((vState = 236) and (hState = 582)) or
								((vState = 236) and (hState = 583)) or
								((vState = 236) and (hState = 584)) or
								((vState = 236) and (hState = 585)) or
								((vState = 236) and (hState = 586)) or
								((vState = 236) and (hState = 587)) or
								((vState = 236) and (hState = 588)) or
								((vState = 236) and (hState = 589)) or
								((vState = 237) and (hState = 557)) or
								((vState = 237) and (hState = 558)) or
								((vState = 237) and (hState = 559)) or
								((vState = 237) and (hState = 560)) or
								((vState = 237) and (hState = 561)) or
								((vState = 237) and (hState = 562)) or
								((vState = 237) and (hState = 563)) or
								((vState = 237) and (hState = 564)) or
								((vState = 237) and (hState = 565)) or
								((vState = 237) and (hState = 566)) or
								((vState = 237) and (hState = 567)) or
								((vState = 237) and (hState = 576)) or
								((vState = 237) and (hState = 577)) or
								((vState = 237) and (hState = 578)) or
								((vState = 237) and (hState = 582)) or
								((vState = 237) and (hState = 583)) or
								((vState = 237) and (hState = 587)) or
								((vState = 237) and (hState = 588)) or
								((vState = 237) and (hState = 589)) or
								((vState = 238) and (hState = 557)) or
								((vState = 238) and (hState = 558)) or
								((vState = 238) and (hState = 559)) or
								((vState = 238) and (hState = 581)) or
								((vState = 238) and (hState = 582)) or
								((vState = 238) and (hState = 583)) or
								((vState = 238) and (hState = 589)) or
								((vState = 239) and (hState = 546)) or
								((vState = 239) and (hState = 547)) or
								((vState = 239) and (hState = 548)) or
								((vState = 239) and (hState = 549)) or
								((vState = 239) and (hState = 550)) or
								((vState = 239) and (hState = 557)) or
								((vState = 239) and (hState = 558)) or
								((vState = 239) and (hState = 582)) or
								((vState = 239) and (hState = 583)) or
								((vState = 240) and (hState = 545)) or
								((vState = 240) and (hState = 546)) or
								((vState = 240) and (hState = 547)) or
								((vState = 240) and (hState = 548)) or
								((vState = 240) and (hState = 549)) or
								((vState = 240) and (hState = 557)) or
								((vState = 240) and (hState = 558)) or
								((vState = 240) and (hState = 574)) or
								((vState = 240) and (hState = 582)) or
								((vState = 240) and (hState = 583)) or
								((vState = 240) and (hState = 584)) or
								((vState = 240) and (hState = 590)) or
								((vState = 240) and (hState = 591)) or
								((vState = 241) and (hState = 537)) or
								((vState = 241) and (hState = 538)) or
								((vState = 241) and (hState = 539)) or
								((vState = 241) and (hState = 540)) or
								((vState = 241) and (hState = 541)) or
								((vState = 241) and (hState = 542)) or
								((vState = 241) and (hState = 543)) or
								((vState = 241) and (hState = 557)) or
								((vState = 241) and (hState = 583)) or
								((vState = 241) and (hState = 584)) or
								((vState = 241) and (hState = 590)) or
								((vState = 241) and (hState = 594)) or
								((vState = 242) and (hState = 531)) or
								((vState = 242) and (hState = 532)) or
								((vState = 242) and (hState = 533)) or
								((vState = 242) and (hState = 534)) or
								((vState = 242) and (hState = 535)) or
								((vState = 242) and (hState = 573)) or
								((vState = 242) and (hState = 584)) or
								((vState = 242) and (hState = 585)) or
								((vState = 242) and (hState = 590)) or
								((vState = 243) and (hState = 556)) or
								((vState = 243) and (hState = 573)) or
								((vState = 243) and (hState = 585)) or
								((vState = 243) and (hState = 586)) or
								((vState = 243) and (hState = 590)) or
								((vState = 244) and (hState = 530)) or
								((vState = 244) and (hState = 587)) or
								((vState = 245) and (hState = 530)) or
								((vState = 245) and (hState = 572)) or
								((vState = 245) and (hState = 588)) or
								((vState = 246) and (hState = 349)) or
								((vState = 246) and (hState = 350)) or
								((vState = 246) and (hState = 530)) or
								((vState = 246) and (hState = 553)) or
								((vState = 246) and (hState = 572)) or
								((vState = 246) and (hState = 588)) or
								((vState = 247) and (hState = 347)) or
								((vState = 247) and (hState = 348)) or
								((vState = 247) and (hState = 349)) or
								((vState = 247) and (hState = 350)) or
								((vState = 247) and (hState = 530)) or
								((vState = 247) and (hState = 542)) or
								((vState = 247) and (hState = 552)) or
								((vState = 247) and (hState = 589)) or
								((vState = 247) and (hState = 590)) or
								((vState = 247) and (hState = 591)) or
								((vState = 248) and (hState = 345)) or
								((vState = 248) and (hState = 346)) or
								((vState = 248) and (hState = 347)) or
								((vState = 248) and (hState = 348)) or
								((vState = 248) and (hState = 530)) or
								((vState = 248) and (hState = 542)) or
								((vState = 249) and (hState = 332)) or
								((vState = 249) and (hState = 347)) or
								((vState = 249) and (hState = 530)) or
								((vState = 249) and (hState = 542)) or
								((vState = 251) and (hState = 323)) or
								((vState = 251) and (hState = 324)) or
								((vState = 251) and (hState = 325)) or
								((vState = 251) and (hState = 335)) or
								((vState = 251) and (hState = 341)) or
								((vState = 251) and (hState = 563)) or
								((vState = 251) and (hState = 569)) or
								((vState = 251) and (hState = 593)) or
								((vState = 252) and (hState = 317)) or
								((vState = 252) and (hState = 318)) or
								((vState = 252) and (hState = 319)) or
								((vState = 252) and (hState = 320)) or
								((vState = 252) and (hState = 321)) or
								((vState = 252) and (hState = 338)) or
								((vState = 252) and (hState = 339)) or
								((vState = 252) and (hState = 340)) or
								((vState = 252) and (hState = 346)) or
								((vState = 252) and (hState = 548)) or
								((vState = 252) and (hState = 563)) or
								((vState = 252) and (hState = 569)) or
								((vState = 252) and (hState = 593)) or
								((vState = 253) and (hState = 312)) or
								((vState = 253) and (hState = 313)) or
								((vState = 253) and (hState = 314)) or
								((vState = 253) and (hState = 315)) or
								((vState = 253) and (hState = 316)) or
								((vState = 253) and (hState = 317)) or
								((vState = 253) and (hState = 318)) or
								((vState = 253) and (hState = 338)) or
								((vState = 253) and (hState = 339)) or
								((vState = 253) and (hState = 340)) or
								((vState = 253) and (hState = 345)) or
								((vState = 253) and (hState = 531)) or
								((vState = 253) and (hState = 541)) or
								((vState = 253) and (hState = 547)) or
								((vState = 253) and (hState = 563)) or
								((vState = 253) and (hState = 568)) or
								((vState = 254) and (hState = 315)) or
								((vState = 254) and (hState = 316)) or
								((vState = 254) and (hState = 341)) or
								((vState = 254) and (hState = 343)) or
								((vState = 254) and (hState = 531)) or
								((vState = 254) and (hState = 541)) or
								((vState = 254) and (hState = 563)) or
								((vState = 254) and (hState = 568)) or
								((vState = 254) and (hState = 594)) or
								((vState = 255) and (hState = 334)) or
								((vState = 255) and (hState = 342)) or
								((vState = 255) and (hState = 343)) or
								((vState = 255) and (hState = 368)) or
								((vState = 255) and (hState = 531)) or
								((vState = 255) and (hState = 541)) or
								((vState = 255) and (hState = 594)) or
								((vState = 256) and (hState = 299)) or
								((vState = 256) and (hState = 300)) or
								((vState = 256) and (hState = 301)) or
								((vState = 256) and (hState = 302)) or
								((vState = 256) and (hState = 303)) or
								((vState = 256) and (hState = 325)) or
								((vState = 256) and (hState = 334)) or
								((vState = 256) and (hState = 343)) or
								((vState = 256) and (hState = 368)) or
								((vState = 256) and (hState = 390)) or
								((vState = 256) and (hState = 531)) or
								((vState = 256) and (hState = 541)) or
								((vState = 256) and (hState = 546)) or
								((vState = 256) and (hState = 594)) or
								((vState = 257) and (hState = 298)) or
								((vState = 257) and (hState = 313)) or
								((vState = 257) and (hState = 326)) or
								((vState = 257) and (hState = 331)) or
								((vState = 257) and (hState = 342)) or
								((vState = 257) and (hState = 343)) or
								((vState = 257) and (hState = 344)) or
								((vState = 257) and (hState = 345)) or
								((vState = 257) and (hState = 371)) or
								((vState = 257) and (hState = 391)) or
								((vState = 257) and (hState = 531)) or
								((vState = 257) and (hState = 562)) or
								((vState = 257) and (hState = 567)) or
								((vState = 257) and (hState = 594)) or
								((vState = 258) and (hState = 328)) or
								((vState = 258) and (hState = 329)) or
								((vState = 258) and (hState = 330)) or
								((vState = 258) and (hState = 341)) or
								((vState = 258) and (hState = 347)) or
								((vState = 258) and (hState = 372)) or
								((vState = 258) and (hState = 373)) or
								((vState = 258) and (hState = 391)) or
								((vState = 258) and (hState = 392)) or
								((vState = 258) and (hState = 531)) or
								((vState = 258) and (hState = 545)) or
								((vState = 258) and (hState = 562)) or
								((vState = 258) and (hState = 567)) or
								((vState = 259) and (hState = 293)) or
								((vState = 259) and (hState = 310)) or
								((vState = 259) and (hState = 328)) or
								((vState = 259) and (hState = 329)) or
								((vState = 259) and (hState = 330)) or
								((vState = 259) and (hState = 340)) or
								((vState = 259) and (hState = 350)) or
								((vState = 259) and (hState = 374)) or
								((vState = 259) and (hState = 392)) or
								((vState = 259) and (hState = 393)) or
								((vState = 259) and (hState = 394)) or
								((vState = 259) and (hState = 531)) or
								((vState = 259) and (hState = 540)) or
								((vState = 259) and (hState = 546)) or
								((vState = 259) and (hState = 557)) or
								((vState = 259) and (hState = 558)) or
								((vState = 259) and (hState = 559)) or
								((vState = 259) and (hState = 560)) or
								((vState = 259) and (hState = 561)) or
								((vState = 259) and (hState = 562)) or
								((vState = 259) and (hState = 563)) or
								((vState = 259) and (hState = 564)) or
								((vState = 259) and (hState = 565)) or
								((vState = 259) and (hState = 566)) or
								((vState = 259) and (hState = 567)) or
								((vState = 259) and (hState = 595)) or
								((vState = 260) and (hState = 292)) or
								((vState = 260) and (hState = 309)) or
								((vState = 260) and (hState = 325)) or
								((vState = 260) and (hState = 331)) or
								((vState = 260) and (hState = 351)) or
								((vState = 260) and (hState = 352)) or
								((vState = 260) and (hState = 377)) or
								((vState = 260) and (hState = 394)) or
								((vState = 260) and (hState = 395)) or
								((vState = 260) and (hState = 540)) or
								((vState = 260) and (hState = 557)) or
								((vState = 260) and (hState = 561)) or
								((vState = 260) and (hState = 569)) or
								((vState = 260) and (hState = 570)) or
								((vState = 260) and (hState = 571)) or
								((vState = 260) and (hState = 572)) or
								((vState = 260) and (hState = 573)) or
								((vState = 260) and (hState = 574)) or
								((vState = 260) and (hState = 575)) or
								((vState = 260) and (hState = 576)) or
								((vState = 260) and (hState = 577)) or
								((vState = 260) and (hState = 578)) or
								((vState = 260) and (hState = 595)) or
								((vState = 261) and (hState = 292)) or
								((vState = 261) and (hState = 309)) or
								((vState = 261) and (hState = 325)) or
								((vState = 261) and (hState = 331)) or
								((vState = 261) and (hState = 351)) or
								((vState = 261) and (hState = 352)) or
								((vState = 261) and (hState = 377)) or
								((vState = 261) and (hState = 394)) or
								((vState = 261) and (hState = 395)) or
								((vState = 261) and (hState = 532)) or
								((vState = 261) and (hState = 540)) or
								((vState = 261) and (hState = 557)) or
								((vState = 261) and (hState = 569)) or
								((vState = 261) and (hState = 570)) or
								((vState = 261) and (hState = 571)) or
								((vState = 261) and (hState = 572)) or
								((vState = 261) and (hState = 573)) or
								((vState = 261) and (hState = 574)) or
								((vState = 261) and (hState = 575)) or
								((vState = 261) and (hState = 576)) or
								((vState = 261) and (hState = 577)) or
								((vState = 261) and (hState = 578)) or
								((vState = 261) and (hState = 595)) or
								((vState = 262) and (hState = 289)) or
								((vState = 262) and (hState = 308)) or
								((vState = 262) and (hState = 324)) or
								((vState = 262) and (hState = 334)) or
								((vState = 262) and (hState = 355)) or
								((vState = 262) and (hState = 378)) or
								((vState = 262) and (hState = 379)) or
								((vState = 262) and (hState = 395)) or
								((vState = 262) and (hState = 396)) or
								((vState = 262) and (hState = 532)) or
								((vState = 262) and (hState = 540)) or
								((vState = 262) and (hState = 550)) or
								((vState = 262) and (hState = 557)) or
								((vState = 262) and (hState = 582)) or
								((vState = 262) and (hState = 583)) or
								((vState = 262) and (hState = 584)) or
								((vState = 262) and (hState = 595)) or
								((vState = 263) and (hState = 287)) or
								((vState = 263) and (hState = 335)) or
								((vState = 263) and (hState = 336)) or
								((vState = 263) and (hState = 337)) or
								((vState = 263) and (hState = 338)) or
								((vState = 263) and (hState = 357)) or
								((vState = 263) and (hState = 358)) or
								((vState = 263) and (hState = 381)) or
								((vState = 263) and (hState = 382)) or
								((vState = 263) and (hState = 396)) or
								((vState = 263) and (hState = 397)) or
								((vState = 263) and (hState = 532)) or
								((vState = 263) and (hState = 551)) or
								((vState = 263) and (hState = 557)) or
								((vState = 263) and (hState = 561)) or
								((vState = 263) and (hState = 588)) or
								((vState = 263) and (hState = 589)) or
								((vState = 263) and (hState = 590)) or
								((vState = 263) and (hState = 591)) or
								((vState = 264) and (hState = 277)) or
								((vState = 264) and (hState = 278)) or
								((vState = 264) and (hState = 279)) or
								((vState = 264) and (hState = 280)) or
								((vState = 264) and (hState = 281)) or
								((vState = 264) and (hState = 282)) or
								((vState = 264) and (hState = 283)) or
								((vState = 264) and (hState = 284)) or
								((vState = 264) and (hState = 285)) or
								((vState = 264) and (hState = 286)) or
								((vState = 264) and (hState = 287)) or
								((vState = 264) and (hState = 304)) or
								((vState = 264) and (hState = 320)) or
								((vState = 264) and (hState = 336)) or
								((vState = 264) and (hState = 337)) or
								((vState = 264) and (hState = 338)) or
								((vState = 264) and (hState = 360)) or
								((vState = 264) and (hState = 361)) or
								((vState = 264) and (hState = 383)) or
								((vState = 264) and (hState = 397)) or
								((vState = 264) and (hState = 398)) or
								((vState = 264) and (hState = 532)) or
								((vState = 264) and (hState = 552)) or
								((vState = 264) and (hState = 561)) or
								((vState = 264) and (hState = 562)) or
								((vState = 264) and (hState = 563)) or
								((vState = 264) and (hState = 588)) or
								((vState = 264) and (hState = 589)) or
								((vState = 264) and (hState = 590)) or
								((vState = 264) and (hState = 591)) or
								((vState = 265) and (hState = 281)) or
								((vState = 265) and (hState = 282)) or
								((vState = 265) and (hState = 283)) or
								((vState = 265) and (hState = 287)) or
								((vState = 265) and (hState = 288)) or
								((vState = 265) and (hState = 289)) or
								((vState = 265) and (hState = 290)) or
								((vState = 265) and (hState = 291)) or
								((vState = 265) and (hState = 292)) or
								((vState = 265) and (hState = 293)) or
								((vState = 265) and (hState = 303)) or
								((vState = 265) and (hState = 318)) or
								((vState = 265) and (hState = 341)) or
								((vState = 265) and (hState = 342)) or
								((vState = 265) and (hState = 343)) or
								((vState = 265) and (hState = 363)) or
								((vState = 265) and (hState = 385)) or
								((vState = 265) and (hState = 397)) or
								((vState = 265) and (hState = 398)) or
								((vState = 265) and (hState = 399)) or
								((vState = 265) and (hState = 400)) or
								((vState = 265) and (hState = 532)) or
								((vState = 265) and (hState = 553)) or
								((vState = 265) and (hState = 558)) or
								((vState = 265) and (hState = 559)) or
								((vState = 265) and (hState = 560)) or
								((vState = 265) and (hState = 561)) or
								((vState = 265) and (hState = 562)) or
								((vState = 265) and (hState = 563)) or
								((vState = 265) and (hState = 585)) or
								((vState = 265) and (hState = 586)) or
								((vState = 266) and (hState = 276)) or
								((vState = 266) and (hState = 281)) or
								((vState = 266) and (hState = 295)) or
								((vState = 266) and (hState = 296)) or
								((vState = 266) and (hState = 297)) or
								((vState = 266) and (hState = 298)) or
								((vState = 266) and (hState = 299)) or
								((vState = 266) and (hState = 300)) or
								((vState = 266) and (hState = 301)) or
								((vState = 266) and (hState = 302)) or
								((vState = 266) and (hState = 303)) or
								((vState = 266) and (hState = 315)) or
								((vState = 266) and (hState = 316)) or
								((vState = 266) and (hState = 335)) or
								((vState = 266) and (hState = 346)) or
								((vState = 266) and (hState = 347)) or
								((vState = 266) and (hState = 348)) or
								((vState = 266) and (hState = 365)) or
								((vState = 266) and (hState = 366)) or
								((vState = 266) and (hState = 367)) or
								((vState = 266) and (hState = 386)) or
								((vState = 266) and (hState = 387)) or
								((vState = 266) and (hState = 388)) or
								((vState = 266) and (hState = 399)) or
								((vState = 266) and (hState = 400)) or
								((vState = 266) and (hState = 401)) or
								((vState = 266) and (hState = 532)) or
								((vState = 266) and (hState = 558)) or
								((vState = 266) and (hState = 559)) or
								((vState = 266) and (hState = 560)) or
								((vState = 266) and (hState = 561)) or
								((vState = 266) and (hState = 562)) or
								((vState = 266) and (hState = 582)) or
								((vState = 266) and (hState = 583)) or
								((vState = 267) and (hState = 276)) or
								((vState = 267) and (hState = 299)) or
								((vState = 267) and (hState = 300)) or
								((vState = 267) and (hState = 301)) or
								((vState = 267) and (hState = 315)) or
								((vState = 267) and (hState = 316)) or
								((vState = 267) and (hState = 366)) or
								((vState = 267) and (hState = 367)) or
								((vState = 267) and (hState = 388)) or
								((vState = 267) and (hState = 399)) or
								((vState = 267) and (hState = 400)) or
								((vState = 267) and (hState = 401)) or
								((vState = 267) and (hState = 532)) or
								((vState = 267) and (hState = 558)) or
								((vState = 267) and (hState = 559)) or
								((vState = 267) and (hState = 560)) or
								((vState = 267) and (hState = 561)) or
								((vState = 267) and (hState = 562)) or
								((vState = 268) and (hState = 276)) or
								((vState = 268) and (hState = 299)) or
								((vState = 268) and (hState = 300)) or
								((vState = 268) and (hState = 309)) or
								((vState = 268) and (hState = 310)) or
								((vState = 268) and (hState = 314)) or
								((vState = 268) and (hState = 315)) or
								((vState = 268) and (hState = 316)) or
								((vState = 268) and (hState = 366)) or
								((vState = 268) and (hState = 367)) or
								((vState = 268) and (hState = 368)) or
								((vState = 268) and (hState = 369)) or
								((vState = 268) and (hState = 371)) or
								((vState = 268) and (hState = 372)) or
								((vState = 268) and (hState = 373)) or
								((vState = 268) and (hState = 374)) or
								((vState = 268) and (hState = 389)) or
								((vState = 268) and (hState = 400)) or
								((vState = 268) and (hState = 401)) or
								((vState = 268) and (hState = 402)) or
								((vState = 268) and (hState = 525)) or
								((vState = 268) and (hState = 558)) or
								((vState = 268) and (hState = 559)) or
								((vState = 268) and (hState = 560)) or
								((vState = 268) and (hState = 561)) or
								((vState = 268) and (hState = 562)) or
								((vState = 269) and (hState = 276)) or
								((vState = 269) and (hState = 277)) or
								((vState = 269) and (hState = 299)) or
								((vState = 269) and (hState = 310)) or
								((vState = 269) and (hState = 311)) or
								((vState = 269) and (hState = 312)) or
								((vState = 269) and (hState = 313)) or
								((vState = 269) and (hState = 314)) or
								((vState = 269) and (hState = 315)) or
								((vState = 269) and (hState = 316)) or
								((vState = 269) and (hState = 317)) or
								((vState = 269) and (hState = 318)) or
								((vState = 269) and (hState = 319)) or
								((vState = 269) and (hState = 320)) or
								((vState = 269) and (hState = 356)) or
								((vState = 269) and (hState = 357)) or
								((vState = 269) and (hState = 365)) or
								((vState = 269) and (hState = 366)) or
								((vState = 269) and (hState = 367)) or
								((vState = 269) and (hState = 368)) or
								((vState = 269) and (hState = 372)) or
								((vState = 269) and (hState = 373)) or
								((vState = 269) and (hState = 374)) or
								((vState = 269) and (hState = 390)) or
								((vState = 269) and (hState = 391)) or
								((vState = 269) and (hState = 401)) or
								((vState = 269) and (hState = 402)) or
								((vState = 269) and (hState = 403)) or
								((vState = 269) and (hState = 525)) or
								((vState = 269) and (hState = 526)) or
								((vState = 269) and (hState = 527)) or
								((vState = 269) and (hState = 558)) or
								((vState = 269) and (hState = 559)) or
								((vState = 269) and (hState = 560)) or
								((vState = 269) and (hState = 561)) or
								((vState = 269) and (hState = 574)) or
								((vState = 269) and (hState = 575)) or
								((vState = 270) and (hState = 275)) or
								((vState = 270) and (hState = 276)) or
								((vState = 270) and (hState = 298)) or
								((vState = 270) and (hState = 310)) or
								((vState = 270) and (hState = 315)) or
								((vState = 270) and (hState = 316)) or
								((vState = 270) and (hState = 317)) or
								((vState = 270) and (hState = 318)) or
								((vState = 270) and (hState = 319)) or
								((vState = 270) and (hState = 320)) or
								((vState = 270) and (hState = 356)) or
								((vState = 270) and (hState = 357)) or
								((vState = 270) and (hState = 358)) or
								((vState = 270) and (hState = 359)) or
								((vState = 270) and (hState = 360)) or
								((vState = 270) and (hState = 361)) or
								((vState = 270) and (hState = 362)) or
								((vState = 270) and (hState = 363)) or
								((vState = 270) and (hState = 364)) or
								((vState = 270) and (hState = 365)) or
								((vState = 270) and (hState = 366)) or
								((vState = 270) and (hState = 367)) or
								((vState = 270) and (hState = 374)) or
								((vState = 270) and (hState = 391)) or
								((vState = 270) and (hState = 392)) or
								((vState = 270) and (hState = 393)) or
								((vState = 270) and (hState = 402)) or
								((vState = 270) and (hState = 403)) or
								((vState = 270) and (hState = 404)) or
								((vState = 270) and (hState = 526)) or
								((vState = 270) and (hState = 527)) or
								((vState = 270) and (hState = 528)) or
								((vState = 270) and (hState = 529)) or
								((vState = 270) and (hState = 560)) or
								((vState = 270) and (hState = 571)) or
								((vState = 270) and (hState = 572)) or
								((vState = 271) and (hState = 273)) or
								((vState = 271) and (hState = 274)) or
								((vState = 271) and (hState = 275)) or
								((vState = 271) and (hState = 276)) or
								((vState = 271) and (hState = 297)) or
								((vState = 271) and (hState = 308)) or
								((vState = 271) and (hState = 309)) or
								((vState = 271) and (hState = 310)) or
								((vState = 271) and (hState = 315)) or
								((vState = 271) and (hState = 316)) or
								((vState = 271) and (hState = 317)) or
								((vState = 271) and (hState = 318)) or
								((vState = 271) and (hState = 319)) or
								((vState = 271) and (hState = 320)) or
								((vState = 271) and (hState = 331)) or
								((vState = 271) and (hState = 354)) or
								((vState = 271) and (hState = 355)) or
								((vState = 271) and (hState = 356)) or
								((vState = 271) and (hState = 364)) or
								((vState = 271) and (hState = 365)) or
								((vState = 271) and (hState = 366)) or
								((vState = 271) and (hState = 367)) or
								((vState = 271) and (hState = 375)) or
								((vState = 271) and (hState = 376)) or
								((vState = 271) and (hState = 377)) or
								((vState = 271) and (hState = 378)) or
								((vState = 271) and (hState = 392)) or
								((vState = 271) and (hState = 393)) or
								((vState = 271) and (hState = 394)) or
								((vState = 271) and (hState = 395)) or
								((vState = 271) and (hState = 402)) or
								((vState = 271) and (hState = 403)) or
								((vState = 271) and (hState = 404)) or
								((vState = 271) and (hState = 405)) or
								((vState = 271) and (hState = 406)) or
								((vState = 271) and (hState = 527)) or
								((vState = 271) and (hState = 528)) or
								((vState = 271) and (hState = 529)) or
								((vState = 271) and (hState = 530)) or
								((vState = 271) and (hState = 560)) or
								((vState = 271) and (hState = 567)) or
								((vState = 271) and (hState = 568)) or
								((vState = 272) and (hState = 276)) or
								((vState = 272) and (hState = 308)) or
								((vState = 272) and (hState = 309)) or
								((vState = 272) and (hState = 310)) or
								((vState = 272) and (hState = 374)) or
								((vState = 272) and (hState = 375)) or
								((vState = 272) and (hState = 376)) or
								((vState = 272) and (hState = 394)) or
								((vState = 272) and (hState = 403)) or
								((vState = 272) and (hState = 404)) or
								((vState = 272) and (hState = 405)) or
								((vState = 272) and (hState = 406)) or
								((vState = 272) and (hState = 527)) or
								((vState = 272) and (hState = 528)) or
								((vState = 272) and (hState = 560)) or
								((vState = 272) and (hState = 561)) or
								((vState = 273) and (hState = 276)) or
								((vState = 273) and (hState = 294)) or
								((vState = 273) and (hState = 308)) or
								((vState = 273) and (hState = 309)) or
								((vState = 273) and (hState = 310)) or
								((vState = 273) and (hState = 329)) or
								((vState = 273) and (hState = 374)) or
								((vState = 273) and (hState = 375)) or
								((vState = 273) and (hState = 379)) or
								((vState = 273) and (hState = 380)) or
								((vState = 273) and (hState = 404)) or
								((vState = 273) and (hState = 405)) or
								((vState = 273) and (hState = 406)) or
								((vState = 273) and (hState = 407)) or
								((vState = 273) and (hState = 528)) or
								((vState = 273) and (hState = 533)) or
								((vState = 273) and (hState = 560)) or
								((vState = 273) and (hState = 561)) or
								((vState = 273) and (hState = 564)) or
								((vState = 274) and (hState = 276)) or
								((vState = 274) and (hState = 293)) or
								((vState = 274) and (hState = 308)) or
								((vState = 274) and (hState = 309)) or
								((vState = 274) and (hState = 329)) or
								((vState = 274) and (hState = 375)) or
								((vState = 274) and (hState = 379)) or
								((vState = 274) and (hState = 380)) or
								((vState = 274) and (hState = 381)) or
								((vState = 274) and (hState = 382)) or
								((vState = 274) and (hState = 383)) or
								((vState = 274) and (hState = 400)) or
								((vState = 274) and (hState = 404)) or
								((vState = 274) and (hState = 405)) or
								((vState = 274) and (hState = 406)) or
								((vState = 274) and (hState = 407)) or
								((vState = 274) and (hState = 408)) or
								((vState = 274) and (hState = 528)) or
								((vState = 274) and (hState = 534)) or
								((vState = 274) and (hState = 558)) or
								((vState = 274) and (hState = 559)) or
								((vState = 274) and (hState = 560)) or
								((vState = 274) and (hState = 599)) or
								((vState = 275) and (hState = 267)) or
								((vState = 275) and (hState = 276)) or
								((vState = 275) and (hState = 292)) or
								((vState = 275) and (hState = 306)) or
								((vState = 275) and (hState = 378)) or
								((vState = 275) and (hState = 379)) or
								((vState = 275) and (hState = 380)) or
								((vState = 275) and (hState = 381)) or
								((vState = 275) and (hState = 382)) or
								((vState = 275) and (hState = 383)) or
								((vState = 275) and (hState = 384)) or
								((vState = 275) and (hState = 385)) or
								((vState = 275) and (hState = 386)) or
								((vState = 275) and (hState = 387)) or
								((vState = 275) and (hState = 401)) or
								((vState = 275) and (hState = 402)) or
								((vState = 275) and (hState = 403)) or
								((vState = 275) and (hState = 404)) or
								((vState = 275) and (hState = 405)) or
								((vState = 275) and (hState = 406)) or
								((vState = 275) and (hState = 529)) or
								((vState = 275) and (hState = 534)) or
								((vState = 275) and (hState = 535)) or
								((vState = 275) and (hState = 540)) or
								((vState = 275) and (hState = 555)) or
								((vState = 275) and (hState = 556)) or
								((vState = 275) and (hState = 557)) or
								((vState = 275) and (hState = 558)) or
								((vState = 275) and (hState = 559)) or
								((vState = 275) and (hState = 574)) or
								((vState = 275) and (hState = 599)) or
								((vState = 276) and (hState = 265)) or
								((vState = 276) and (hState = 276)) or
								((vState = 276) and (hState = 302)) or
								((vState = 276) and (hState = 303)) or
								((vState = 276) and (hState = 335)) or
								((vState = 276) and (hState = 336)) or
								((vState = 276) and (hState = 337)) or
								((vState = 276) and (hState = 373)) or
								((vState = 276) and (hState = 383)) or
								((vState = 276) and (hState = 384)) or
								((vState = 276) and (hState = 385)) or
								((vState = 276) and (hState = 386)) or
								((vState = 276) and (hState = 387)) or
								((vState = 276) and (hState = 388)) or
								((vState = 276) and (hState = 389)) or
								((vState = 276) and (hState = 404)) or
								((vState = 276) and (hState = 405)) or
								((vState = 276) and (hState = 406)) or
								((vState = 276) and (hState = 411)) or
								((vState = 276) and (hState = 529)) or
								((vState = 276) and (hState = 534)) or
								((vState = 276) and (hState = 540)) or
								((vState = 276) and (hState = 551)) or
								((vState = 276) and (hState = 552)) or
								((vState = 276) and (hState = 558)) or
								((vState = 276) and (hState = 559)) or
								((vState = 276) and (hState = 567)) or
								((vState = 276) and (hState = 574)) or
								((vState = 276) and (hState = 599)) or
								((vState = 277) and (hState = 276)) or
								((vState = 277) and (hState = 373)) or
								((vState = 277) and (hState = 387)) or
								((vState = 277) and (hState = 388)) or
								((vState = 277) and (hState = 389)) or
								((vState = 277) and (hState = 406)) or
								((vState = 277) and (hState = 540)) or
								((vState = 277) and (hState = 558)) or
								((vState = 277) and (hState = 559)) or
								((vState = 277) and (hState = 560)) or
								((vState = 277) and (hState = 574)) or
								((vState = 278) and (hState = 262)) or
								((vState = 278) and (hState = 276)) or
								((vState = 278) and (hState = 326)) or
								((vState = 278) and (hState = 327)) or
								((vState = 278) and (hState = 373)) or
								((vState = 278) and (hState = 397)) or
								((vState = 278) and (hState = 540)) or
								((vState = 278) and (hState = 558)) or
								((vState = 278) and (hState = 559)) or
								((vState = 278) and (hState = 560)) or
								((vState = 278) and (hState = 574)) or
								((vState = 278) and (hState = 588)) or
								((vState = 279) and (hState = 262)) or
								((vState = 279) and (hState = 276)) or
								((vState = 279) and (hState = 294)) or
								((vState = 279) and (hState = 325)) or
								((vState = 279) and (hState = 326)) or
								((vState = 279) and (hState = 327)) or
								((vState = 279) and (hState = 328)) or
								((vState = 279) and (hState = 340)) or
								((vState = 279) and (hState = 373)) or
								((vState = 279) and (hState = 395)) or
								((vState = 279) and (hState = 396)) or
								((vState = 279) and (hState = 530)) or
								((vState = 279) and (hState = 535)) or
								((vState = 279) and (hState = 540)) or
								((vState = 279) and (hState = 544)) or
								((vState = 279) and (hState = 557)) or
								((vState = 279) and (hState = 558)) or
								((vState = 279) and (hState = 559)) or
								((vState = 279) and (hState = 560)) or
								((vState = 279) and (hState = 574)) or
								((vState = 279) and (hState = 575)) or
								((vState = 279) and (hState = 588)) or
								((vState = 280) and (hState = 262)) or
								((vState = 280) and (hState = 276)) or
								((vState = 280) and (hState = 293)) or
								((vState = 280) and (hState = 325)) or
								((vState = 280) and (hState = 326)) or
								((vState = 280) and (hState = 327)) or
								((vState = 280) and (hState = 341)) or
								((vState = 280) and (hState = 373)) or
								((vState = 280) and (hState = 374)) or
								((vState = 280) and (hState = 375)) or
								((vState = 280) and (hState = 376)) or
								((vState = 280) and (hState = 377)) or
								((vState = 280) and (hState = 378)) or
								((vState = 280) and (hState = 379)) or
								((vState = 280) and (hState = 400)) or
								((vState = 280) and (hState = 535)) or
								((vState = 280) and (hState = 540)) or
								((vState = 280) and (hState = 541)) or
								((vState = 280) and (hState = 542)) or
								((vState = 280) and (hState = 543)) or
								((vState = 280) and (hState = 557)) or
								((vState = 280) and (hState = 558)) or
								((vState = 280) and (hState = 559)) or
								((vState = 280) and (hState = 560)) or
								((vState = 280) and (hState = 572)) or
								((vState = 280) and (hState = 573)) or
								((vState = 280) and (hState = 574)) or
								((vState = 280) and (hState = 575)) or
								((vState = 280) and (hState = 588)) or
								((vState = 281) and (hState = 262)) or
								((vState = 281) and (hState = 276)) or
								((vState = 281) and (hState = 324)) or
								((vState = 281) and (hState = 342)) or
								((vState = 281) and (hState = 368)) or
								((vState = 281) and (hState = 369)) or
								((vState = 281) and (hState = 370)) or
								((vState = 281) and (hState = 371)) or
								((vState = 281) and (hState = 372)) or
								((vState = 281) and (hState = 373)) or
								((vState = 281) and (hState = 401)) or
								((vState = 281) and (hState = 531)) or
								((vState = 281) and (hState = 535)) or
								((vState = 281) and (hState = 536)) or
								((vState = 281) and (hState = 537)) or
								((vState = 281) and (hState = 541)) or
								((vState = 281) and (hState = 542)) or
								((vState = 281) and (hState = 543)) or
								((vState = 281) and (hState = 556)) or
								((vState = 281) and (hState = 557)) or
								((vState = 281) and (hState = 558)) or
								((vState = 281) and (hState = 559)) or
								((vState = 281) and (hState = 560)) or
								((vState = 281) and (hState = 573)) or
								((vState = 281) and (hState = 574)) or
								((vState = 281) and (hState = 575)) or
								((vState = 282) and (hState = 276)) or
								((vState = 282) and (hState = 323)) or
								((vState = 282) and (hState = 324)) or
								((vState = 282) and (hState = 343)) or
								((vState = 282) and (hState = 402)) or
								((vState = 282) and (hState = 531)) or
								((vState = 282) and (hState = 532)) or
								((vState = 282) and (hState = 535)) or
								((vState = 282) and (hState = 541)) or
								((vState = 282) and (hState = 556)) or
								((vState = 282) and (hState = 560)) or
								((vState = 282) and (hState = 574)) or
								((vState = 282) and (hState = 575)) or
								((vState = 282) and (hState = 576)) or
								((vState = 283) and (hState = 276)) or
								((vState = 283) and (hState = 320)) or
								((vState = 283) and (hState = 321)) or
								((vState = 283) and (hState = 322)) or
								((vState = 283) and (hState = 323)) or
								((vState = 283) and (hState = 324)) or
								((vState = 283) and (hState = 342)) or
								((vState = 283) and (hState = 343)) or
								((vState = 283) and (hState = 362)) or
								((vState = 283) and (hState = 367)) or
								((vState = 283) and (hState = 531)) or
								((vState = 283) and (hState = 532)) or
								((vState = 283) and (hState = 533)) or
								((vState = 283) and (hState = 534)) or
								((vState = 283) and (hState = 535)) or
								((vState = 283) and (hState = 560)) or
								((vState = 283) and (hState = 561)) or
								((vState = 283) and (hState = 575)) or
								((vState = 283) and (hState = 576)) or
								((vState = 283) and (hState = 577)) or
								((vState = 283) and (hState = 589)) or
								((vState = 284) and (hState = 276)) or
								((vState = 284) and (hState = 310)) or
								((vState = 284) and (hState = 311)) or
								((vState = 284) and (hState = 312)) or
								((vState = 284) and (hState = 313)) or
								((vState = 284) and (hState = 314)) or
								((vState = 284) and (hState = 315)) or
								((vState = 284) and (hState = 316)) or
								((vState = 284) and (hState = 317)) or
								((vState = 284) and (hState = 344)) or
								((vState = 284) and (hState = 345)) or
								((vState = 284) and (hState = 346)) or
								((vState = 284) and (hState = 347)) or
								((vState = 284) and (hState = 348)) or
								((vState = 284) and (hState = 349)) or
								((vState = 284) and (hState = 350)) or
								((vState = 284) and (hState = 351)) or
								((vState = 284) and (hState = 352)) or
								((vState = 284) and (hState = 353)) or
								((vState = 284) and (hState = 354)) or
								((vState = 284) and (hState = 355)) or
								((vState = 284) and (hState = 531)) or
								((vState = 284) and (hState = 532)) or
								((vState = 284) and (hState = 533)) or
								((vState = 284) and (hState = 534)) or
								((vState = 284) and (hState = 535)) or
								((vState = 284) and (hState = 560)) or
								((vState = 284) and (hState = 561)) or
								((vState = 284) and (hState = 562)) or
								((vState = 284) and (hState = 576)) or
								((vState = 284) and (hState = 577)) or
								((vState = 284) and (hState = 589)) or
								((vState = 285) and (hState = 276)) or
								((vState = 285) and (hState = 281)) or
								((vState = 285) and (hState = 309)) or
								((vState = 285) and (hState = 310)) or
								((vState = 285) and (hState = 311)) or
								((vState = 285) and (hState = 312)) or
								((vState = 285) and (hState = 313)) or
								((vState = 285) and (hState = 314)) or
								((vState = 285) and (hState = 315)) or
								((vState = 285) and (hState = 316)) or
								((vState = 285) and (hState = 345)) or
								((vState = 285) and (hState = 346)) or
								((vState = 285) and (hState = 347)) or
								((vState = 285) and (hState = 348)) or
								((vState = 285) and (hState = 349)) or
								((vState = 285) and (hState = 350)) or
								((vState = 285) and (hState = 351)) or
								((vState = 285) and (hState = 352)) or
								((vState = 285) and (hState = 353)) or
								((vState = 285) and (hState = 354)) or
								((vState = 285) and (hState = 355)) or
								((vState = 285) and (hState = 370)) or
								((vState = 285) and (hState = 371)) or
								((vState = 285) and (hState = 372)) or
								((vState = 285) and (hState = 405)) or
								((vState = 285) and (hState = 531)) or
								((vState = 285) and (hState = 532)) or
								((vState = 285) and (hState = 533)) or
								((vState = 285) and (hState = 534)) or
								((vState = 285) and (hState = 535)) or
								((vState = 285) and (hState = 542)) or
								((vState = 285) and (hState = 548)) or
								((vState = 285) and (hState = 560)) or
								((vState = 285) and (hState = 561)) or
								((vState = 285) and (hState = 562)) or
								((vState = 285) and (hState = 576)) or
								((vState = 285) and (hState = 577)) or
								((vState = 285) and (hState = 578)) or
								((vState = 285) and (hState = 589)) or
								((vState = 286) and (hState = 276)) or
								((vState = 286) and (hState = 281)) or
								((vState = 286) and (hState = 289)) or
								((vState = 286) and (hState = 309)) or
								((vState = 286) and (hState = 310)) or
								((vState = 286) and (hState = 311)) or
								((vState = 286) and (hState = 312)) or
								((vState = 286) and (hState = 313)) or
								((vState = 286) and (hState = 345)) or
								((vState = 286) and (hState = 346)) or
								((vState = 286) and (hState = 347)) or
								((vState = 286) and (hState = 348)) or
								((vState = 286) and (hState = 372)) or
								((vState = 286) and (hState = 406)) or
								((vState = 286) and (hState = 531)) or
								((vState = 286) and (hState = 532)) or
								((vState = 286) and (hState = 533)) or
								((vState = 286) and (hState = 534)) or
								((vState = 286) and (hState = 535)) or
								((vState = 286) and (hState = 542)) or
								((vState = 286) and (hState = 560)) or
								((vState = 286) and (hState = 561)) or
								((vState = 286) and (hState = 562)) or
								((vState = 286) and (hState = 576)) or
								((vState = 286) and (hState = 577)) or
								((vState = 286) and (hState = 578)) or
								((vState = 286) and (hState = 579)) or
								((vState = 286) and (hState = 590)) or
								((vState = 287) and (hState = 276)) or
								((vState = 287) and (hState = 281)) or
								((vState = 287) and (hState = 288)) or
								((vState = 287) and (hState = 306)) or
								((vState = 287) and (hState = 307)) or
								((vState = 287) and (hState = 308)) or
								((vState = 287) and (hState = 309)) or
								((vState = 287) and (hState = 310)) or
								((vState = 287) and (hState = 338)) or
								((vState = 287) and (hState = 339)) or
								((vState = 287) and (hState = 340)) or
								((vState = 287) and (hState = 341)) or
								((vState = 287) and (hState = 342)) or
								((vState = 287) and (hState = 343)) or
								((vState = 287) and (hState = 344)) or
								((vState = 287) and (hState = 345)) or
								((vState = 287) and (hState = 346)) or
								((vState = 287) and (hState = 347)) or
								((vState = 287) and (hState = 348)) or
								((vState = 287) and (hState = 372)) or
								((vState = 287) and (hState = 373)) or
								((vState = 287) and (hState = 374)) or
								((vState = 287) and (hState = 407)) or
								((vState = 287) and (hState = 531)) or
								((vState = 287) and (hState = 532)) or
								((vState = 287) and (hState = 535)) or
								((vState = 287) and (hState = 542)) or
								((vState = 287) and (hState = 552)) or
								((vState = 287) and (hState = 553)) or
								((vState = 287) and (hState = 561)) or
								((vState = 287) and (hState = 562)) or
								((vState = 287) and (hState = 579)) or
								((vState = 287) and (hState = 580)) or
								((vState = 287) and (hState = 590)) or
								((vState = 288) and (hState = 276)) or
								((vState = 288) and (hState = 288)) or
								((vState = 288) and (hState = 305)) or
								((vState = 288) and (hState = 306)) or
								((vState = 288) and (hState = 307)) or
								((vState = 288) and (hState = 308)) or
								((vState = 288) and (hState = 340)) or
								((vState = 288) and (hState = 341)) or
								((vState = 288) and (hState = 342)) or
								((vState = 288) and (hState = 372)) or
								((vState = 288) and (hState = 535)) or
								((vState = 288) and (hState = 552)) or
								((vState = 288) and (hState = 553)) or
								((vState = 288) and (hState = 561)) or
								((vState = 288) and (hState = 562)) or
								((vState = 288) and (hState = 579)) or
								((vState = 288) and (hState = 580)) or
								((vState = 288) and (hState = 590)) or
								((vState = 289) and (hState = 276)) or
								((vState = 289) and (hState = 302)) or
								((vState = 289) and (hState = 303)) or
								((vState = 289) and (hState = 304)) or
								((vState = 289) and (hState = 305)) or
								((vState = 289) and (hState = 306)) or
								((vState = 289) and (hState = 336)) or
								((vState = 289) and (hState = 340)) or
								((vState = 289) and (hState = 350)) or
								((vState = 289) and (hState = 372)) or
								((vState = 289) and (hState = 536)) or
								((vState = 289) and (hState = 552)) or
								((vState = 289) and (hState = 553)) or
								((vState = 289) and (hState = 561)) or
								((vState = 289) and (hState = 562)) or
								((vState = 289) and (hState = 579)) or
								((vState = 289) and (hState = 580)) or
								((vState = 289) and (hState = 581)) or
								((vState = 290) and (hState = 276)) or
								((vState = 290) and (hState = 287)) or
								((vState = 290) and (hState = 298)) or
								((vState = 290) and (hState = 299)) or
								((vState = 290) and (hState = 300)) or
								((vState = 290) and (hState = 301)) or
								((vState = 290) and (hState = 302)) or
								((vState = 290) and (hState = 303)) or
								((vState = 290) and (hState = 304)) or
								((vState = 290) and (hState = 305)) or
								((vState = 290) and (hState = 336)) or
								((vState = 290) and (hState = 340)) or
								((vState = 290) and (hState = 351)) or
								((vState = 290) and (hState = 372)) or
								((vState = 290) and (hState = 378)) or
								((vState = 290) and (hState = 423)) or
								((vState = 290) and (hState = 532)) or
								((vState = 290) and (hState = 536)) or
								((vState = 290) and (hState = 552)) or
								((vState = 290) and (hState = 553)) or
								((vState = 290) and (hState = 554)) or
								((vState = 290) and (hState = 561)) or
								((vState = 290) and (hState = 562)) or
								((vState = 290) and (hState = 563)) or
								((vState = 290) and (hState = 577)) or
								((vState = 290) and (hState = 578)) or
								((vState = 290) and (hState = 579)) or
								((vState = 290) and (hState = 580)) or
								((vState = 290) and (hState = 581)) or
								((vState = 290) and (hState = 582)) or
								((vState = 290) and (hState = 583)) or
								((vState = 291) and (hState = 276)) or
								((vState = 291) and (hState = 294)) or
								((vState = 291) and (hState = 295)) or
								((vState = 291) and (hState = 296)) or
								((vState = 291) and (hState = 297)) or
								((vState = 291) and (hState = 298)) or
								((vState = 291) and (hState = 299)) or
								((vState = 291) and (hState = 300)) or
								((vState = 291) and (hState = 301)) or
								((vState = 291) and (hState = 335)) or
								((vState = 291) and (hState = 336)) or
								((vState = 291) and (hState = 337)) or
								((vState = 291) and (hState = 352)) or
								((vState = 291) and (hState = 378)) or
								((vState = 291) and (hState = 379)) or
								((vState = 291) and (hState = 380)) or
								((vState = 291) and (hState = 532)) or
								((vState = 291) and (hState = 536)) or
								((vState = 291) and (hState = 557)) or
								((vState = 291) and (hState = 562)) or
								((vState = 291) and (hState = 563)) or
								((vState = 291) and (hState = 577)) or
								((vState = 291) and (hState = 581)) or
								((vState = 291) and (hState = 582)) or
								((vState = 291) and (hState = 583)) or
								((vState = 291) and (hState = 584)) or
								((vState = 292) and (hState = 294)) or
								((vState = 292) and (hState = 295)) or
								((vState = 292) and (hState = 296)) or
								((vState = 292) and (hState = 297)) or
								((vState = 292) and (hState = 298)) or
								((vState = 292) and (hState = 299)) or
								((vState = 292) and (hState = 335)) or
								((vState = 292) and (hState = 353)) or
								((vState = 292) and (hState = 371)) or
								((vState = 292) and (hState = 375)) or
								((vState = 292) and (hState = 376)) or
								((vState = 292) and (hState = 377)) or
								((vState = 292) and (hState = 378)) or
								((vState = 292) and (hState = 381)) or
								((vState = 292) and (hState = 382)) or
								((vState = 292) and (hState = 388)) or
								((vState = 292) and (hState = 389)) or
								((vState = 292) and (hState = 390)) or
								((vState = 292) and (hState = 391)) or
								((vState = 292) and (hState = 392)) or
								((vState = 292) and (hState = 532)) or
								((vState = 292) and (hState = 536)) or
								((vState = 292) and (hState = 551)) or
								((vState = 292) and (hState = 558)) or
								((vState = 292) and (hState = 562)) or
								((vState = 292) and (hState = 563)) or
								((vState = 292) and (hState = 577)) or
								((vState = 292) and (hState = 583)) or
								((vState = 292) and (hState = 584)) or
								((vState = 292) and (hState = 585)) or
								((vState = 292) and (hState = 586)) or
								((vState = 293) and (hState = 294)) or
								((vState = 293) and (hState = 295)) or
								((vState = 293) and (hState = 335)) or
								((vState = 293) and (hState = 370)) or
								((vState = 293) and (hState = 371)) or
								((vState = 293) and (hState = 374)) or
								((vState = 293) and (hState = 375)) or
								((vState = 293) and (hState = 376)) or
								((vState = 293) and (hState = 377)) or
								((vState = 293) and (hState = 378)) or
								((vState = 293) and (hState = 382)) or
								((vState = 293) and (hState = 536)) or
								((vState = 293) and (hState = 551)) or
								((vState = 293) and (hState = 562)) or
								((vState = 293) and (hState = 563)) or
								((vState = 293) and (hState = 577)) or
								((vState = 293) and (hState = 584)) or
								((vState = 293) and (hState = 585)) or
								((vState = 293) and (hState = 586)) or
								((vState = 293) and (hState = 587)) or
								((vState = 294) and (hState = 266)) or
								((vState = 294) and (hState = 293)) or
								((vState = 294) and (hState = 333)) or
								((vState = 294) and (hState = 334)) or
								((vState = 294) and (hState = 335)) or
								((vState = 294) and (hState = 354)) or
								((vState = 294) and (hState = 355)) or
								((vState = 294) and (hState = 369)) or
								((vState = 294) and (hState = 370)) or
								((vState = 294) and (hState = 371)) or
								((vState = 294) and (hState = 372)) or
								((vState = 294) and (hState = 373)) or
								((vState = 294) and (hState = 374)) or
								((vState = 294) and (hState = 375)) or
								((vState = 294) and (hState = 376)) or
								((vState = 294) and (hState = 377)) or
								((vState = 294) and (hState = 378)) or
								((vState = 294) and (hState = 386)) or
								((vState = 294) and (hState = 387)) or
								((vState = 294) and (hState = 405)) or
								((vState = 294) and (hState = 406)) or
								((vState = 294) and (hState = 536)) or
								((vState = 294) and (hState = 537)) or
								((vState = 294) and (hState = 562)) or
								((vState = 294) and (hState = 563)) or
								((vState = 294) and (hState = 577)) or
								((vState = 294) and (hState = 585)) or
								((vState = 294) and (hState = 586)) or
								((vState = 294) and (hState = 587)) or
								((vState = 294) and (hState = 588)) or
								((vState = 295) and (hState = 266)) or
								((vState = 295) and (hState = 278)) or
								((vState = 295) and (hState = 293)) or
								((vState = 295) and (hState = 325)) or
								((vState = 295) and (hState = 326)) or
								((vState = 295) and (hState = 327)) or
								((vState = 295) and (hState = 328)) or
								((vState = 295) and (hState = 329)) or
								((vState = 295) and (hState = 330)) or
								((vState = 295) and (hState = 331)) or
								((vState = 295) and (hState = 332)) or
								((vState = 295) and (hState = 333)) or
								((vState = 295) and (hState = 334)) or
								((vState = 295) and (hState = 335)) or
								((vState = 295) and (hState = 336)) or
								((vState = 295) and (hState = 337)) or
								((vState = 295) and (hState = 338)) or
								((vState = 295) and (hState = 339)) or
								((vState = 295) and (hState = 340)) or
								((vState = 295) and (hState = 341)) or
								((vState = 295) and (hState = 342)) or
								((vState = 295) and (hState = 343)) or
								((vState = 295) and (hState = 344)) or
								((vState = 295) and (hState = 345)) or
								((vState = 295) and (hState = 346)) or
								((vState = 295) and (hState = 347)) or
								((vState = 295) and (hState = 348)) or
								((vState = 295) and (hState = 349)) or
								((vState = 295) and (hState = 350)) or
								((vState = 295) and (hState = 351)) or
								((vState = 295) and (hState = 352)) or
								((vState = 295) and (hState = 353)) or
								((vState = 295) and (hState = 354)) or
								((vState = 295) and (hState = 355)) or
								((vState = 295) and (hState = 356)) or
								((vState = 295) and (hState = 357)) or
								((vState = 295) and (hState = 358)) or
								((vState = 295) and (hState = 363)) or
								((vState = 295) and (hState = 364)) or
								((vState = 295) and (hState = 365)) or
								((vState = 295) and (hState = 366)) or
								((vState = 295) and (hState = 370)) or
								((vState = 295) and (hState = 371)) or
								((vState = 295) and (hState = 372)) or
								((vState = 295) and (hState = 373)) or
								((vState = 295) and (hState = 374)) or
								((vState = 295) and (hState = 375)) or
								((vState = 295) and (hState = 376)) or
								((vState = 295) and (hState = 377)) or
								((vState = 295) and (hState = 378)) or
								((vState = 295) and (hState = 386)) or
								((vState = 295) and (hState = 387)) or
								((vState = 295) and (hState = 395)) or
								((vState = 295) and (hState = 405)) or
								((vState = 295) and (hState = 406)) or
								((vState = 295) and (hState = 413)) or
								((vState = 295) and (hState = 428)) or
								((vState = 295) and (hState = 534)) or
								((vState = 295) and (hState = 535)) or
								((vState = 295) and (hState = 536)) or
								((vState = 295) and (hState = 537)) or
								((vState = 295) and (hState = 562)) or
								((vState = 295) and (hState = 563)) or
								((vState = 295) and (hState = 564)) or
								((vState = 295) and (hState = 577)) or
								((vState = 295) and (hState = 585)) or
								((vState = 295) and (hState = 586)) or
								((vState = 295) and (hState = 587)) or
								((vState = 295) and (hState = 588)) or
								((vState = 295) and (hState = 589)) or
								((vState = 295) and (hState = 590)) or
								((vState = 295) and (hState = 591)) or
								((vState = 296) and (hState = 266)) or
								((vState = 296) and (hState = 278)) or
								((vState = 296) and (hState = 283)) or
								((vState = 296) and (hState = 289)) or
								((vState = 296) and (hState = 290)) or
								((vState = 296) and (hState = 291)) or
								((vState = 296) and (hState = 292)) or
								((vState = 296) and (hState = 293)) or
								((vState = 296) and (hState = 320)) or
								((vState = 296) and (hState = 325)) or
								((vState = 296) and (hState = 326)) or
								((vState = 296) and (hState = 327)) or
								((vState = 296) and (hState = 357)) or
								((vState = 296) and (hState = 358)) or
								((vState = 296) and (hState = 362)) or
								((vState = 296) and (hState = 363)) or
								((vState = 296) and (hState = 364)) or
								((vState = 296) and (hState = 365)) or
								((vState = 296) and (hState = 366)) or
								((vState = 296) and (hState = 370)) or
								((vState = 296) and (hState = 371)) or
								((vState = 296) and (hState = 372)) or
								((vState = 296) and (hState = 388)) or
								((vState = 296) and (hState = 389)) or
								((vState = 296) and (hState = 397)) or
								((vState = 296) and (hState = 405)) or
								((vState = 296) and (hState = 406)) or
								((vState = 296) and (hState = 429)) or
								((vState = 296) and (hState = 534)) or
								((vState = 296) and (hState = 535)) or
								((vState = 296) and (hState = 536)) or
								((vState = 296) and (hState = 537)) or
								((vState = 296) and (hState = 538)) or
								((vState = 296) and (hState = 563)) or
								((vState = 296) and (hState = 564)) or
								((vState = 296) and (hState = 588)) or
								((vState = 296) and (hState = 589)) or
								((vState = 296) and (hState = 590)) or
								((vState = 296) and (hState = 591)) or
								((vState = 297) and (hState = 278)) or
								((vState = 297) and (hState = 282)) or
								((vState = 297) and (hState = 283)) or
								((vState = 297) and (hState = 287)) or
								((vState = 297) and (hState = 288)) or
								((vState = 297) and (hState = 293)) or
								((vState = 297) and (hState = 320)) or
								((vState = 297) and (hState = 324)) or
								((vState = 297) and (hState = 325)) or
								((vState = 297) and (hState = 357)) or
								((vState = 297) and (hState = 358)) or
								((vState = 297) and (hState = 362)) or
								((vState = 297) and (hState = 363)) or
								((vState = 297) and (hState = 364)) or
								((vState = 297) and (hState = 365)) or
								((vState = 297) and (hState = 366)) or
								((vState = 297) and (hState = 367)) or
								((vState = 297) and (hState = 371)) or
								((vState = 297) and (hState = 390)) or
								((vState = 297) and (hState = 404)) or
								((vState = 297) and (hState = 405)) or
								((vState = 297) and (hState = 406)) or
								((vState = 297) and (hState = 416)) or
								((vState = 297) and (hState = 534)) or
								((vState = 297) and (hState = 535)) or
								((vState = 297) and (hState = 548)) or
								((vState = 297) and (hState = 563)) or
								((vState = 297) and (hState = 564)) or
								((vState = 297) and (hState = 565)) or
								((vState = 297) and (hState = 578)) or
								((vState = 297) and (hState = 589)) or
								((vState = 297) and (hState = 590)) or
								((vState = 297) and (hState = 591)) or
								((vState = 298) and (hState = 282)) or
								((vState = 298) and (hState = 283)) or
								((vState = 298) and (hState = 293)) or
								((vState = 298) and (hState = 320)) or
								((vState = 298) and (hState = 357)) or
								((vState = 298) and (hState = 358)) or
								((vState = 298) and (hState = 362)) or
								((vState = 298) and (hState = 363)) or
								((vState = 298) and (hState = 364)) or
								((vState = 298) and (hState = 371)) or
								((vState = 298) and (hState = 404)) or
								((vState = 298) and (hState = 405)) or
								((vState = 298) and (hState = 406)) or
								((vState = 298) and (hState = 534)) or
								((vState = 298) and (hState = 535)) or
								((vState = 298) and (hState = 548)) or
								((vState = 298) and (hState = 563)) or
								((vState = 298) and (hState = 564)) or
								((vState = 298) and (hState = 565)) or
								((vState = 298) and (hState = 566)) or
								((vState = 298) and (hState = 578)) or
								((vState = 298) and (hState = 590)) or
								((vState = 298) and (hState = 591)) or
								((vState = 298) and (hState = 592)) or
								((vState = 299) and (hState = 267)) or
								((vState = 299) and (hState = 282)) or
								((vState = 299) and (hState = 293)) or
								((vState = 299) and (hState = 319)) or
								((vState = 299) and (hState = 320)) or
								((vState = 299) and (hState = 357)) or
								((vState = 299) and (hState = 358)) or
								((vState = 299) and (hState = 359)) or
								((vState = 299) and (hState = 360)) or
								((vState = 299) and (hState = 361)) or
								((vState = 299) and (hState = 362)) or
								((vState = 299) and (hState = 406)) or
								((vState = 299) and (hState = 534)) or
								((vState = 299) and (hState = 535)) or
								((vState = 299) and (hState = 540)) or
								((vState = 299) and (hState = 546)) or
								((vState = 299) and (hState = 564)) or
								((vState = 299) and (hState = 565)) or
								((vState = 299) and (hState = 566)) or
								((vState = 299) and (hState = 567)) or
								((vState = 299) and (hState = 578)) or
								((vState = 299) and (hState = 593)) or
								((vState = 300) and (hState = 275)) or
								((vState = 300) and (hState = 276)) or
								((vState = 300) and (hState = 277)) or
								((vState = 300) and (hState = 293)) or
								((vState = 300) and (hState = 351)) or
								((vState = 300) and (hState = 352)) or
								((vState = 300) and (hState = 353)) or
								((vState = 300) and (hState = 354)) or
								((vState = 300) and (hState = 355)) or
								((vState = 300) and (hState = 356)) or
								((vState = 300) and (hState = 357)) or
								((vState = 300) and (hState = 358)) or
								((vState = 300) and (hState = 359)) or
								((vState = 300) and (hState = 360)) or
								((vState = 300) and (hState = 361)) or
								((vState = 300) and (hState = 362)) or
								((vState = 300) and (hState = 402)) or
								((vState = 300) and (hState = 418)) or
								((vState = 300) and (hState = 530)) or
								((vState = 300) and (hState = 531)) or
								((vState = 300) and (hState = 532)) or
								((vState = 300) and (hState = 533)) or
								((vState = 300) and (hState = 534)) or
								((vState = 300) and (hState = 535)) or
								((vState = 300) and (hState = 540)) or
								((vState = 300) and (hState = 546)) or
								((vState = 300) and (hState = 565)) or
								((vState = 300) and (hState = 566)) or
								((vState = 300) and (hState = 578)) or
								((vState = 300) and (hState = 595)) or
								((vState = 301) and (hState = 275)) or
								((vState = 301) and (hState = 276)) or
								((vState = 301) and (hState = 277)) or
								((vState = 301) and (hState = 293)) or
								((vState = 301) and (hState = 330)) or
								((vState = 301) and (hState = 351)) or
								((vState = 301) and (hState = 352)) or
								((vState = 301) and (hState = 353)) or
								((vState = 301) and (hState = 354)) or
								((vState = 301) and (hState = 355)) or
								((vState = 301) and (hState = 356)) or
								((vState = 301) and (hState = 357)) or
								((vState = 301) and (hState = 358)) or
								((vState = 301) and (hState = 359)) or
								((vState = 301) and (hState = 360)) or
								((vState = 301) and (hState = 361)) or
								((vState = 301) and (hState = 362)) or
								((vState = 301) and (hState = 396)) or
								((vState = 301) and (hState = 402)) or
								((vState = 301) and (hState = 418)) or
								((vState = 301) and (hState = 434)) or
								((vState = 301) and (hState = 518)) or
								((vState = 301) and (hState = 519)) or
								((vState = 301) and (hState = 530)) or
								((vState = 301) and (hState = 531)) or
								((vState = 301) and (hState = 532)) or
								((vState = 301) and (hState = 533)) or
								((vState = 301) and (hState = 534)) or
								((vState = 301) and (hState = 535)) or
								((vState = 301) and (hState = 540)) or
								((vState = 301) and (hState = 541)) or
								((vState = 301) and (hState = 546)) or
								((vState = 301) and (hState = 565)) or
								((vState = 301) and (hState = 578)) or
								((vState = 301) and (hState = 589)) or
								((vState = 301) and (hState = 595)) or
								((vState = 301) and (hState = 596)) or
								((vState = 302) and (hState = 275)) or
								((vState = 302) and (hState = 276)) or
								((vState = 302) and (hState = 277)) or
								((vState = 302) and (hState = 293)) or
								((vState = 302) and (hState = 314)) or
								((vState = 302) and (hState = 315)) or
								((vState = 302) and (hState = 354)) or
								((vState = 302) and (hState = 355)) or
								((vState = 302) and (hState = 356)) or
								((vState = 302) and (hState = 357)) or
								((vState = 302) and (hState = 363)) or
								((vState = 302) and (hState = 364)) or
								((vState = 302) and (hState = 365)) or
								((vState = 302) and (hState = 366)) or
								((vState = 302) and (hState = 367)) or
								((vState = 302) and (hState = 368)) or
								((vState = 302) and (hState = 369)) or
								((vState = 302) and (hState = 370)) or
								((vState = 302) and (hState = 371)) or
								((vState = 302) and (hState = 372)) or
								((vState = 302) and (hState = 402)) or
								((vState = 302) and (hState = 403)) or
								((vState = 302) and (hState = 407)) or
								((vState = 302) and (hState = 418)) or
								((vState = 302) and (hState = 517)) or
								((vState = 302) and (hState = 530)) or
								((vState = 302) and (hState = 535)) or
								((vState = 302) and (hState = 536)) or
								((vState = 302) and (hState = 537)) or
								((vState = 302) and (hState = 538)) or
								((vState = 302) and (hState = 539)) or
								((vState = 302) and (hState = 540)) or
								((vState = 302) and (hState = 541)) or
								((vState = 302) and (hState = 545)) or
								((vState = 302) and (hState = 546)) or
								((vState = 302) and (hState = 565)) or
								((vState = 302) and (hState = 571)) or
								((vState = 302) and (hState = 572)) or
								((vState = 302) and (hState = 578)) or
								((vState = 302) and (hState = 597)) or
								((vState = 303) and (hState = 275)) or
								((vState = 303) and (hState = 276)) or
								((vState = 303) and (hState = 293)) or
								((vState = 303) and (hState = 313)) or
								((vState = 303) and (hState = 314)) or
								((vState = 303) and (hState = 329)) or
								((vState = 303) and (hState = 354)) or
								((vState = 303) and (hState = 355)) or
								((vState = 303) and (hState = 364)) or
								((vState = 303) and (hState = 369)) or
								((vState = 303) and (hState = 402)) or
								((vState = 303) and (hState = 403)) or
								((vState = 303) and (hState = 404)) or
								((vState = 303) and (hState = 406)) or
								((vState = 303) and (hState = 407)) or
								((vState = 303) and (hState = 418)) or
								((vState = 303) and (hState = 529)) or
								((vState = 303) and (hState = 536)) or
								((vState = 303) and (hState = 541)) or
								((vState = 303) and (hState = 542)) or
								((vState = 303) and (hState = 544)) or
								((vState = 303) and (hState = 545)) or
								((vState = 303) and (hState = 546)) or
								((vState = 303) and (hState = 547)) or
								((vState = 303) and (hState = 564)) or
								((vState = 303) and (hState = 565)) or
								((vState = 303) and (hState = 566)) or
								((vState = 303) and (hState = 573)) or
								((vState = 303) and (hState = 588)) or
								((vState = 303) and (hState = 598)) or
								((vState = 304) and (hState = 275)) or
								((vState = 304) and (hState = 276)) or
								((vState = 304) and (hState = 293)) or
								((vState = 304) and (hState = 313)) or
								((vState = 304) and (hState = 384)) or
								((vState = 304) and (hState = 401)) or
								((vState = 304) and (hState = 402)) or
								((vState = 304) and (hState = 403)) or
								((vState = 304) and (hState = 404)) or
								((vState = 304) and (hState = 405)) or
								((vState = 304) and (hState = 406)) or
								((vState = 304) and (hState = 407)) or
								((vState = 304) and (hState = 418)) or
								((vState = 304) and (hState = 536)) or
								((vState = 304) and (hState = 542)) or
								((vState = 304) and (hState = 543)) or
								((vState = 304) and (hState = 544)) or
								((vState = 304) and (hState = 545)) or
								((vState = 304) and (hState = 546)) or
								((vState = 304) and (hState = 547)) or
								((vState = 305) and (hState = 275)) or
								((vState = 305) and (hState = 276)) or
								((vState = 305) and (hState = 293)) or
								((vState = 305) and (hState = 304)) or
								((vState = 305) and (hState = 384)) or
								((vState = 305) and (hState = 385)) or
								((vState = 305) and (hState = 386)) or
								((vState = 305) and (hState = 387)) or
								((vState = 305) and (hState = 388)) or
								((vState = 305) and (hState = 401)) or
								((vState = 305) and (hState = 402)) or
								((vState = 305) and (hState = 403)) or
								((vState = 305) and (hState = 404)) or
								((vState = 305) and (hState = 405)) or
								((vState = 305) and (hState = 406)) or
								((vState = 305) and (hState = 407)) or
								((vState = 305) and (hState = 536)) or
								((vState = 305) and (hState = 542)) or
								((vState = 305) and (hState = 543)) or
								((vState = 305) and (hState = 544)) or
								((vState = 305) and (hState = 547)) or
								((vState = 305) and (hState = 556)) or
								((vState = 306) and (hState = 275)) or
								((vState = 306) and (hState = 276)) or
								((vState = 306) and (hState = 293)) or
								((vState = 306) and (hState = 304)) or
								((vState = 306) and (hState = 305)) or
								((vState = 306) and (hState = 306)) or
								((vState = 306) and (hState = 335)) or
								((vState = 306) and (hState = 336)) or
								((vState = 306) and (hState = 337)) or
								((vState = 306) and (hState = 338)) or
								((vState = 306) and (hState = 339)) or
								((vState = 306) and (hState = 340)) or
								((vState = 306) and (hState = 349)) or
								((vState = 306) and (hState = 350)) or
								((vState = 306) and (hState = 384)) or
								((vState = 306) and (hState = 385)) or
								((vState = 306) and (hState = 386)) or
								((vState = 306) and (hState = 387)) or
								((vState = 306) and (hState = 388)) or
								((vState = 306) and (hState = 399)) or
								((vState = 306) and (hState = 400)) or
								((vState = 306) and (hState = 401)) or
								((vState = 306) and (hState = 402)) or
								((vState = 306) and (hState = 403)) or
								((vState = 306) and (hState = 404)) or
								((vState = 306) and (hState = 405)) or
								((vState = 306) and (hState = 406)) or
								((vState = 306) and (hState = 407)) or
								((vState = 306) and (hState = 408)) or
								((vState = 306) and (hState = 432)) or
								((vState = 306) and (hState = 433)) or
								((vState = 306) and (hState = 439)) or
								((vState = 306) and (hState = 511)) or
								((vState = 306) and (hState = 526)) or
								((vState = 306) and (hState = 527)) or
								((vState = 306) and (hState = 536)) or
								((vState = 306) and (hState = 542)) or
								((vState = 306) and (hState = 543)) or
								((vState = 306) and (hState = 547)) or
								((vState = 306) and (hState = 548)) or
								((vState = 306) and (hState = 549)) or
								((vState = 306) and (hState = 550)) or
								((vState = 306) and (hState = 551)) or
								((vState = 306) and (hState = 552)) or
								((vState = 306) and (hState = 553)) or
								((vState = 306) and (hState = 554)) or
								((vState = 306) and (hState = 555)) or
								((vState = 306) and (hState = 556)) or
								((vState = 306) and (hState = 577)) or
								((vState = 307) and (hState = 275)) or
								((vState = 307) and (hState = 276)) or
								((vState = 307) and (hState = 303)) or
								((vState = 307) and (hState = 304)) or
								((vState = 307) and (hState = 342)) or
								((vState = 307) and (hState = 343)) or
								((vState = 307) and (hState = 344)) or
								((vState = 307) and (hState = 345)) or
								((vState = 307) and (hState = 346)) or
								((vState = 307) and (hState = 347)) or
								((vState = 307) and (hState = 348)) or
								((vState = 307) and (hState = 349)) or
								((vState = 307) and (hState = 350)) or
								((vState = 307) and (hState = 368)) or
								((vState = 307) and (hState = 388)) or
								((vState = 307) and (hState = 400)) or
								((vState = 307) and (hState = 401)) or
								((vState = 307) and (hState = 402)) or
								((vState = 307) and (hState = 403)) or
								((vState = 307) and (hState = 404)) or
								((vState = 307) and (hState = 405)) or
								((vState = 307) and (hState = 406)) or
								((vState = 307) and (hState = 407)) or
								((vState = 307) and (hState = 408)) or
								((vState = 307) and (hState = 409)) or
								((vState = 307) and (hState = 417)) or
								((vState = 307) and (hState = 429)) or
								((vState = 307) and (hState = 434)) or
								((vState = 307) and (hState = 508)) or
								((vState = 307) and (hState = 525)) or
								((vState = 307) and (hState = 536)) or
								((vState = 307) and (hState = 541)) or
								((vState = 307) and (hState = 542)) or
								((vState = 307) and (hState = 543)) or
								((vState = 307) and (hState = 547)) or
								((vState = 307) and (hState = 548)) or
								((vState = 307) and (hState = 549)) or
								((vState = 307) and (hState = 553)) or
								((vState = 307) and (hState = 554)) or
								((vState = 307) and (hState = 555)) or
								((vState = 307) and (hState = 556)) or
								((vState = 307) and (hState = 566)) or
								((vState = 307) and (hState = 567)) or
								((vState = 307) and (hState = 579)) or
								((vState = 308) and (hState = 301)) or
								((vState = 308) and (hState = 302)) or
								((vState = 308) and (hState = 303)) or
								((vState = 308) and (hState = 304)) or
								((vState = 308) and (hState = 310)) or
								((vState = 308) and (hState = 311)) or
								((vState = 308) and (hState = 326)) or
								((vState = 308) and (hState = 334)) or
								((vState = 308) and (hState = 343)) or
								((vState = 308) and (hState = 344)) or
								((vState = 308) and (hState = 345)) or
								((vState = 308) and (hState = 346)) or
								((vState = 308) and (hState = 347)) or
								((vState = 308) and (hState = 348)) or
								((vState = 308) and (hState = 349)) or
								((vState = 308) and (hState = 350)) or
								((vState = 308) and (hState = 351)) or
								((vState = 308) and (hState = 361)) or
								((vState = 308) and (hState = 368)) or
								((vState = 308) and (hState = 383)) or
								((vState = 308) and (hState = 390)) or
								((vState = 308) and (hState = 400)) or
								((vState = 308) and (hState = 406)) or
								((vState = 308) and (hState = 407)) or
								((vState = 308) and (hState = 408)) or
								((vState = 308) and (hState = 409)) or
								((vState = 308) and (hState = 410)) or
								((vState = 308) and (hState = 411)) or
								((vState = 308) and (hState = 417)) or
								((vState = 308) and (hState = 427)) or
								((vState = 308) and (hState = 507)) or
								((vState = 308) and (hState = 524)) or
								((vState = 308) and (hState = 536)) or
								((vState = 308) and (hState = 540)) or
								((vState = 308) and (hState = 541)) or
								((vState = 308) and (hState = 542)) or
								((vState = 308) and (hState = 543)) or
								((vState = 308) and (hState = 544)) or
								((vState = 308) and (hState = 545)) or
								((vState = 308) and (hState = 548)) or
								((vState = 308) and (hState = 558)) or
								((vState = 308) and (hState = 559)) or
								((vState = 308) and (hState = 566)) or
								((vState = 308) and (hState = 567)) or
								((vState = 308) and (hState = 585)) or
								((vState = 309) and (hState = 304)) or
								((vState = 309) and (hState = 310)) or
								((vState = 309) and (hState = 311)) or
								((vState = 309) and (hState = 361)) or
								((vState = 309) and (hState = 368)) or
								((vState = 309) and (hState = 400)) or
								((vState = 309) and (hState = 408)) or
								((vState = 309) and (hState = 409)) or
								((vState = 309) and (hState = 410)) or
								((vState = 309) and (hState = 411)) or
								((vState = 309) and (hState = 417)) or
								((vState = 309) and (hState = 536)) or
								((vState = 309) and (hState = 540)) or
								((vState = 309) and (hState = 541)) or
								((vState = 309) and (hState = 566)) or
								((vState = 309) and (hState = 567)) or
								((vState = 310) and (hState = 299)) or
								((vState = 310) and (hState = 304)) or
								((vState = 310) and (hState = 309)) or
								((vState = 310) and (hState = 310)) or
								((vState = 310) and (hState = 361)) or
								((vState = 310) and (hState = 368)) or
								((vState = 310) and (hState = 382)) or
								((vState = 310) and (hState = 409)) or
								((vState = 310) and (hState = 412)) or
								((vState = 310) and (hState = 413)) or
								((vState = 310) and (hState = 417)) or
								((vState = 310) and (hState = 536)) or
								((vState = 310) and (hState = 537)) or
								((vState = 310) and (hState = 538)) or
								((vState = 310) and (hState = 539)) or
								((vState = 310) and (hState = 540)) or
								((vState = 310) and (hState = 567)) or
								((vState = 311) and (hState = 292)) or
								((vState = 311) and (hState = 299)) or
								((vState = 311) and (hState = 304)) or
								((vState = 311) and (hState = 308)) or
								((vState = 311) and (hState = 309)) or
								((vState = 311) and (hState = 310)) or
								((vState = 311) and (hState = 325)) or
								((vState = 311) and (hState = 331)) or
								((vState = 311) and (hState = 359)) or
								((vState = 311) and (hState = 360)) or
								((vState = 311) and (hState = 361)) or
								((vState = 311) and (hState = 362)) or
								((vState = 311) and (hState = 368)) or
								((vState = 311) and (hState = 381)) or
								((vState = 311) and (hState = 382)) or
								((vState = 311) and (hState = 394)) or
								((vState = 311) and (hState = 395)) or
								((vState = 311) and (hState = 412)) or
								((vState = 311) and (hState = 413)) or
								((vState = 311) and (hState = 414)) or
								((vState = 311) and (hState = 415)) or
								((vState = 311) and (hState = 416)) or
								((vState = 311) and (hState = 417)) or
								((vState = 311) and (hState = 423)) or
								((vState = 311) and (hState = 438)) or
								((vState = 311) and (hState = 444)) or
								((vState = 311) and (hState = 502)) or
								((vState = 311) and (hState = 503)) or
								((vState = 311) and (hState = 522)) or
								((vState = 311) and (hState = 530)) or
								((vState = 311) and (hState = 531)) or
								((vState = 311) and (hState = 532)) or
								((vState = 311) and (hState = 533)) or
								((vState = 311) and (hState = 534)) or
								((vState = 311) and (hState = 535)) or
								((vState = 311) and (hState = 536)) or
								((vState = 311) and (hState = 537)) or
								((vState = 311) and (hState = 538)) or
								((vState = 311) and (hState = 539)) or
								((vState = 311) and (hState = 540)) or
								((vState = 311) and (hState = 567)) or
								((vState = 311) and (hState = 568)) or
								((vState = 311) and (hState = 584)) or
								((vState = 312) and (hState = 271)) or
								((vState = 312) and (hState = 292)) or
								((vState = 312) and (hState = 299)) or
								((vState = 312) and (hState = 304)) or
								((vState = 312) and (hState = 308)) or
								((vState = 312) and (hState = 309)) or
								((vState = 312) and (hState = 310)) or
								((vState = 312) and (hState = 336)) or
								((vState = 312) and (hState = 359)) or
								((vState = 312) and (hState = 360)) or
								((vState = 312) and (hState = 361)) or
								((vState = 312) and (hState = 365)) or
								((vState = 312) and (hState = 366)) or
								((vState = 312) and (hState = 367)) or
								((vState = 312) and (hState = 368)) or
								((vState = 312) and (hState = 372)) or
								((vState = 312) and (hState = 396)) or
								((vState = 312) and (hState = 397)) or
								((vState = 312) and (hState = 398)) or
								((vState = 312) and (hState = 415)) or
								((vState = 312) and (hState = 416)) or
								((vState = 312) and (hState = 417)) or
								((vState = 312) and (hState = 421)) or
								((vState = 312) and (hState = 439)) or
								((vState = 312) and (hState = 501)) or
								((vState = 312) and (hState = 529)) or
								((vState = 312) and (hState = 530)) or
								((vState = 312) and (hState = 531)) or
								((vState = 312) and (hState = 536)) or
								((vState = 312) and (hState = 537)) or
								((vState = 312) and (hState = 538)) or
								((vState = 312) and (hState = 539)) or
								((vState = 312) and (hState = 540)) or
								((vState = 312) and (hState = 567)) or
								((vState = 312) and (hState = 568)) or
								((vState = 312) and (hState = 569)) or
								((vState = 312) and (hState = 570)) or
								((vState = 312) and (hState = 571)) or
								((vState = 312) and (hState = 572)) or
								((vState = 312) and (hState = 573)) or
								((vState = 312) and (hState = 584)) or
								((vState = 312) and (hState = 585)) or
								((vState = 313) and (hState = 271)) or
								((vState = 313) and (hState = 292)) or
								((vState = 313) and (hState = 299)) or
								((vState = 313) and (hState = 304)) or
								((vState = 313) and (hState = 305)) or
								((vState = 313) and (hState = 306)) or
								((vState = 313) and (hState = 307)) or
								((vState = 313) and (hState = 308)) or
								((vState = 313) and (hState = 309)) or
								((vState = 313) and (hState = 310)) or
								((vState = 313) and (hState = 324)) or
								((vState = 313) and (hState = 330)) or
								((vState = 313) and (hState = 334)) or
								((vState = 313) and (hState = 361)) or
								((vState = 313) and (hState = 368)) or
								((vState = 313) and (hState = 369)) or
								((vState = 313) and (hState = 370)) or
								((vState = 313) and (hState = 371)) or
								((vState = 313) and (hState = 372)) or
								((vState = 313) and (hState = 373)) or
								((vState = 313) and (hState = 416)) or
								((vState = 313) and (hState = 417)) or
								((vState = 313) and (hState = 418)) or
								((vState = 313) and (hState = 419)) or
								((vState = 313) and (hState = 420)) or
								((vState = 313) and (hState = 421)) or
								((vState = 313) and (hState = 519)) or
								((vState = 313) and (hState = 525)) or
								((vState = 313) and (hState = 526)) or
								((vState = 313) and (hState = 527)) or
								((vState = 313) and (hState = 528)) or
								((vState = 313) and (hState = 536)) or
								((vState = 313) and (hState = 537)) or
								((vState = 313) and (hState = 538)) or
								((vState = 313) and (hState = 539)) or
								((vState = 313) and (hState = 540)) or
								((vState = 313) and (hState = 541)) or
								((vState = 313) and (hState = 568)) or
								((vState = 313) and (hState = 576)) or
								((vState = 313) and (hState = 577)) or
								((vState = 313) and (hState = 583)) or
								((vState = 314) and (hState = 271)) or
								((vState = 314) and (hState = 292)) or
								((vState = 314) and (hState = 299)) or
								((vState = 314) and (hState = 304)) or
								((vState = 314) and (hState = 305)) or
								((vState = 314) and (hState = 306)) or
								((vState = 314) and (hState = 307)) or
								((vState = 314) and (hState = 308)) or
								((vState = 314) and (hState = 309)) or
								((vState = 314) and (hState = 330)) or
								((vState = 314) and (hState = 361)) or
								((vState = 314) and (hState = 368)) or
								((vState = 314) and (hState = 416)) or
								((vState = 314) and (hState = 417)) or
								((vState = 314) and (hState = 519)) or
								((vState = 314) and (hState = 526)) or
								((vState = 314) and (hState = 527)) or
								((vState = 314) and (hState = 528)) or
								((vState = 314) and (hState = 539)) or
								((vState = 314) and (hState = 568)) or
								((vState = 314) and (hState = 583)) or
								((vState = 315) and (hState = 272)) or
								((vState = 315) and (hState = 273)) or
								((vState = 315) and (hState = 274)) or
								((vState = 315) and (hState = 292)) or
								((vState = 315) and (hState = 299)) or
								((vState = 315) and (hState = 304)) or
								((vState = 315) and (hState = 305)) or
								((vState = 315) and (hState = 309)) or
								((vState = 315) and (hState = 329)) or
								((vState = 315) and (hState = 357)) or
								((vState = 315) and (hState = 361)) or
								((vState = 315) and (hState = 368)) or
								((vState = 315) and (hState = 375)) or
								((vState = 315) and (hState = 376)) or
								((vState = 315) and (hState = 377)) or
								((vState = 315) and (hState = 378)) or
								((vState = 315) and (hState = 379)) or
								((vState = 315) and (hState = 416)) or
								((vState = 315) and (hState = 518)) or
								((vState = 315) and (hState = 527)) or
								((vState = 315) and (hState = 535)) or
								((vState = 315) and (hState = 568)) or
								((vState = 316) and (hState = 272)) or
								((vState = 316) and (hState = 273)) or
								((vState = 316) and (hState = 274)) or
								((vState = 316) and (hState = 292)) or
								((vState = 316) and (hState = 299)) or
								((vState = 316) and (hState = 304)) or
								((vState = 316) and (hState = 305)) or
								((vState = 316) and (hState = 309)) or
								((vState = 316) and (hState = 328)) or
								((vState = 316) and (hState = 349)) or
								((vState = 316) and (hState = 350)) or
								((vState = 316) and (hState = 353)) or
								((vState = 316) and (hState = 354)) or
								((vState = 316) and (hState = 355)) or
								((vState = 316) and (hState = 356)) or
								((vState = 316) and (hState = 359)) or
								((vState = 316) and (hState = 360)) or
								((vState = 316) and (hState = 361)) or
								((vState = 316) and (hState = 368)) or
								((vState = 316) and (hState = 376)) or
								((vState = 316) and (hState = 377)) or
								((vState = 316) and (hState = 378)) or
								((vState = 316) and (hState = 379)) or
								((vState = 316) and (hState = 380)) or
								((vState = 316) and (hState = 381)) or
								((vState = 316) and (hState = 382)) or
								((vState = 316) and (hState = 383)) or
								((vState = 316) and (hState = 384)) or
								((vState = 316) and (hState = 397)) or
								((vState = 316) and (hState = 403)) or
								((vState = 316) and (hState = 415)) or
								((vState = 316) and (hState = 416)) or
								((vState = 316) and (hState = 443)) or
								((vState = 316) and (hState = 449)) or
								((vState = 316) and (hState = 516)) or
								((vState = 316) and (hState = 518)) or
								((vState = 316) and (hState = 526)) or
								((vState = 316) and (hState = 534)) or
								((vState = 316) and (hState = 535)) or
								((vState = 316) and (hState = 549)) or
								((vState = 316) and (hState = 568)) or
								((vState = 317) and (hState = 272)) or
								((vState = 317) and (hState = 273)) or
								((vState = 317) and (hState = 274)) or
								((vState = 317) and (hState = 292)) or
								((vState = 317) and (hState = 303)) or
								((vState = 317) and (hState = 304)) or
								((vState = 317) and (hState = 309)) or
								((vState = 317) and (hState = 323)) or
								((vState = 317) and (hState = 324)) or
								((vState = 317) and (hState = 325)) or
								((vState = 317) and (hState = 326)) or
								((vState = 317) and (hState = 355)) or
								((vState = 317) and (hState = 361)) or
								((vState = 317) and (hState = 362)) or
								((vState = 317) and (hState = 363)) or
								((vState = 317) and (hState = 364)) or
								((vState = 317) and (hState = 365)) or
								((vState = 317) and (hState = 366)) or
								((vState = 317) and (hState = 367)) or
								((vState = 317) and (hState = 368)) or
								((vState = 317) and (hState = 369)) or
								((vState = 317) and (hState = 370)) or
								((vState = 317) and (hState = 371)) or
								((vState = 317) and (hState = 376)) or
								((vState = 317) and (hState = 377)) or
								((vState = 317) and (hState = 378)) or
								((vState = 317) and (hState = 379)) or
								((vState = 317) and (hState = 380)) or
								((vState = 317) and (hState = 381)) or
								((vState = 317) and (hState = 382)) or
								((vState = 317) and (hState = 383)) or
								((vState = 317) and (hState = 386)) or
								((vState = 317) and (hState = 387)) or
								((vState = 317) and (hState = 388)) or
								((vState = 317) and (hState = 389)) or
								((vState = 317) and (hState = 397)) or
								((vState = 317) and (hState = 405)) or
								((vState = 317) and (hState = 413)) or
								((vState = 317) and (hState = 414)) or
								((vState = 317) and (hState = 415)) or
								((vState = 317) and (hState = 416)) or
								((vState = 317) and (hState = 428)) or
								((vState = 317) and (hState = 429)) or
								((vState = 317) and (hState = 444)) or
								((vState = 317) and (hState = 492)) or
								((vState = 317) and (hState = 493)) or
								((vState = 317) and (hState = 512)) or
								((vState = 317) and (hState = 513)) or
								((vState = 317) and (hState = 514)) or
								((vState = 317) and (hState = 525)) or
								((vState = 317) and (hState = 531)) or
								((vState = 317) and (hState = 532)) or
								((vState = 317) and (hState = 533)) or
								((vState = 317) and (hState = 534)) or
								((vState = 317) and (hState = 551)) or
								((vState = 317) and (hState = 552)) or
								((vState = 317) and (hState = 553)) or
								((vState = 317) and (hState = 568)) or
								((vState = 317) and (hState = 593)) or
								((vState = 318) and (hState = 272)) or
								((vState = 318) and (hState = 273)) or
								((vState = 318) and (hState = 274)) or
								((vState = 318) and (hState = 292)) or
								((vState = 318) and (hState = 302)) or
								((vState = 318) and (hState = 303)) or
								((vState = 318) and (hState = 304)) or
								((vState = 318) and (hState = 308)) or
								((vState = 318) and (hState = 322)) or
								((vState = 318) and (hState = 323)) or
								((vState = 318) and (hState = 324)) or
								((vState = 318) and (hState = 325)) or
								((vState = 318) and (hState = 326)) or
								((vState = 318) and (hState = 347)) or
								((vState = 318) and (hState = 355)) or
								((vState = 318) and (hState = 361)) or
								((vState = 318) and (hState = 367)) or
								((vState = 318) and (hState = 374)) or
								((vState = 318) and (hState = 375)) or
								((vState = 318) and (hState = 376)) or
								((vState = 318) and (hState = 377)) or
								((vState = 318) and (hState = 378)) or
								((vState = 318) and (hState = 379)) or
								((vState = 318) and (hState = 380)) or
								((vState = 318) and (hState = 381)) or
								((vState = 318) and (hState = 382)) or
								((vState = 318) and (hState = 383)) or
								((vState = 318) and (hState = 391)) or
								((vState = 318) and (hState = 392)) or
								((vState = 318) and (hState = 393)) or
								((vState = 318) and (hState = 394)) or
								((vState = 318) and (hState = 395)) or
								((vState = 318) and (hState = 396)) or
								((vState = 318) and (hState = 397)) or
								((vState = 318) and (hState = 407)) or
								((vState = 318) and (hState = 408)) or
								((vState = 318) and (hState = 409)) or
								((vState = 318) and (hState = 410)) or
								((vState = 318) and (hState = 411)) or
								((vState = 318) and (hState = 491)) or
								((vState = 318) and (hState = 507)) or
								((vState = 318) and (hState = 508)) or
								((vState = 318) and (hState = 509)) or
								((vState = 318) and (hState = 510)) or
								((vState = 318) and (hState = 511)) or
								((vState = 318) and (hState = 512)) or
								((vState = 318) and (hState = 513)) or
								((vState = 318) and (hState = 524)) or
								((vState = 318) and (hState = 530)) or
								((vState = 318) and (hState = 531)) or
								((vState = 318) and (hState = 532)) or
								((vState = 318) and (hState = 533)) or
								((vState = 318) and (hState = 551)) or
								((vState = 318) and (hState = 556)) or
								((vState = 318) and (hState = 557)) or
								((vState = 318) and (hState = 594)) or
								((vState = 319) and (hState = 272)) or
								((vState = 319) and (hState = 273)) or
								((vState = 319) and (hState = 274)) or
								((vState = 319) and (hState = 292)) or
								((vState = 319) and (hState = 302)) or
								((vState = 319) and (hState = 303)) or
								((vState = 319) and (hState = 304)) or
								((vState = 319) and (hState = 308)) or
								((vState = 319) and (hState = 321)) or
								((vState = 319) and (hState = 322)) or
								((vState = 319) and (hState = 323)) or
								((vState = 319) and (hState = 324)) or
								((vState = 319) and (hState = 325)) or
								((vState = 319) and (hState = 347)) or
								((vState = 319) and (hState = 361)) or
								((vState = 319) and (hState = 367)) or
								((vState = 319) and (hState = 375)) or
								((vState = 319) and (hState = 379)) or
								((vState = 319) and (hState = 380)) or
								((vState = 319) and (hState = 396)) or
								((vState = 319) and (hState = 397)) or
								((vState = 319) and (hState = 407)) or
								((vState = 319) and (hState = 408)) or
								((vState = 319) and (hState = 409)) or
								((vState = 319) and (hState = 410)) or
								((vState = 319) and (hState = 411)) or
								((vState = 319) and (hState = 511)) or
								((vState = 319) and (hState = 512)) or
								((vState = 319) and (hState = 530)) or
								((vState = 319) and (hState = 531)) or
								((vState = 319) and (hState = 532)) or
								((vState = 319) and (hState = 551)) or
								((vState = 320) and (hState = 272)) or
								((vState = 320) and (hState = 273)) or
								((vState = 320) and (hState = 274)) or
								((vState = 320) and (hState = 292)) or
								((vState = 320) and (hState = 298)) or
								((vState = 320) and (hState = 320)) or
								((vState = 320) and (hState = 321)) or
								((vState = 320) and (hState = 322)) or
								((vState = 320) and (hState = 323)) or
								((vState = 320) and (hState = 324)) or
								((vState = 320) and (hState = 325)) or
								((vState = 320) and (hState = 361)) or
								((vState = 320) and (hState = 367)) or
								((vState = 320) and (hState = 380)) or
								((vState = 320) and (hState = 396)) or
								((vState = 320) and (hState = 407)) or
								((vState = 320) and (hState = 408)) or
								((vState = 320) and (hState = 409)) or
								((vState = 320) and (hState = 410)) or
								((vState = 320) and (hState = 411)) or
								((vState = 320) and (hState = 511)) or
								((vState = 320) and (hState = 521)) or
								((vState = 320) and (hState = 522)) or
								((vState = 320) and (hState = 523)) or
								((vState = 320) and (hState = 530)) or
								((vState = 320) and (hState = 531)) or
								((vState = 320) and (hState = 532)) or
								((vState = 320) and (hState = 551)) or
								((vState = 321) and (hState = 272)) or
								((vState = 321) and (hState = 273)) or
								((vState = 321) and (hState = 274)) or
								((vState = 321) and (hState = 292)) or
								((vState = 321) and (hState = 298)) or
								((vState = 321) and (hState = 299)) or
								((vState = 321) and (hState = 300)) or
								((vState = 321) and (hState = 322)) or
								((vState = 321) and (hState = 323)) or
								((vState = 321) and (hState = 324)) or
								((vState = 321) and (hState = 325)) or
								((vState = 321) and (hState = 361)) or
								((vState = 321) and (hState = 367)) or
								((vState = 321) and (hState = 410)) or
								((vState = 321) and (hState = 413)) or
								((vState = 321) and (hState = 414)) or
								((vState = 321) and (hState = 522)) or
								((vState = 321) and (hState = 523)) or
								((vState = 321) and (hState = 526)) or
								((vState = 321) and (hState = 527)) or
								((vState = 321) and (hState = 530)) or
								((vState = 321) and (hState = 540)) or
								((vState = 322) and (hState = 272)) or
								((vState = 322) and (hState = 273)) or
								((vState = 322) and (hState = 274)) or
								((vState = 322) and (hState = 292)) or
								((vState = 322) and (hState = 298)) or
								((vState = 322) and (hState = 299)) or
								((vState = 322) and (hState = 323)) or
								((vState = 322) and (hState = 324)) or
								((vState = 322) and (hState = 325)) or
								((vState = 322) and (hState = 346)) or
								((vState = 322) and (hState = 352)) or
								((vState = 322) and (hState = 361)) or
								((vState = 322) and (hState = 367)) or
								((vState = 322) and (hState = 382)) or
								((vState = 322) and (hState = 395)) or
								((vState = 322) and (hState = 402)) or
								((vState = 322) and (hState = 403)) or
								((vState = 322) and (hState = 404)) or
								((vState = 322) and (hState = 405)) or
								((vState = 322) and (hState = 406)) or
								((vState = 322) and (hState = 413)) or
								((vState = 322) and (hState = 414)) or
								((vState = 322) and (hState = 454)) or
								((vState = 322) and (hState = 485)) or
								((vState = 322) and (hState = 503)) or
								((vState = 322) and (hState = 522)) or
								((vState = 322) and (hState = 523)) or
								((vState = 322) and (hState = 524)) or
								((vState = 322) and (hState = 525)) or
								((vState = 322) and (hState = 526)) or
								((vState = 322) and (hState = 527)) or
								((vState = 322) and (hState = 530)) or
								((vState = 322) and (hState = 540)) or
								((vState = 322) and (hState = 567)) or
								((vState = 322) and (hState = 568)) or
								((vState = 322) and (hState = 569)) or
								((vState = 322) and (hState = 599)) or
								((vState = 323) and (hState = 272)) or
								((vState = 323) and (hState = 273)) or
								((vState = 323) and (hState = 292)) or
								((vState = 323) and (hState = 298)) or
								((vState = 323) and (hState = 299)) or
								((vState = 323) and (hState = 304)) or
								((vState = 323) and (hState = 305)) or
								((vState = 323) and (hState = 306)) or
								((vState = 323) and (hState = 319)) or
								((vState = 323) and (hState = 328)) or
								((vState = 323) and (hState = 329)) or
								((vState = 323) and (hState = 351)) or
								((vState = 323) and (hState = 361)) or
								((vState = 323) and (hState = 367)) or
								((vState = 323) and (hState = 383)) or
								((vState = 323) and (hState = 395)) or
								((vState = 323) and (hState = 402)) or
								((vState = 323) and (hState = 403)) or
								((vState = 323) and (hState = 404)) or
								((vState = 323) and (hState = 405)) or
								((vState = 323) and (hState = 406)) or
								((vState = 323) and (hState = 415)) or
								((vState = 323) and (hState = 416)) or
								((vState = 323) and (hState = 455)) or
								((vState = 323) and (hState = 483)) or
								((vState = 323) and (hState = 508)) or
								((vState = 323) and (hState = 521)) or
								((vState = 323) and (hState = 522)) or
								((vState = 323) and (hState = 523)) or
								((vState = 323) and (hState = 528)) or
								((vState = 323) and (hState = 529)) or
								((vState = 323) and (hState = 530)) or
								((vState = 323) and (hState = 540)) or
								((vState = 323) and (hState = 552)) or
								((vState = 323) and (hState = 571)) or
								((vState = 323) and (hState = 572)) or
								((vState = 323) and (hState = 573)) or
								((vState = 324) and (hState = 271)) or
								((vState = 324) and (hState = 272)) or
								((vState = 324) and (hState = 273)) or
								((vState = 324) and (hState = 292)) or
								((vState = 324) and (hState = 297)) or
								((vState = 324) and (hState = 298)) or
								((vState = 324) and (hState = 304)) or
								((vState = 324) and (hState = 305)) or
								((vState = 324) and (hState = 319)) or
								((vState = 324) and (hState = 320)) or
								((vState = 324) and (hState = 321)) or
								((vState = 324) and (hState = 331)) or
								((vState = 324) and (hState = 332)) or
								((vState = 324) and (hState = 345)) or
								((vState = 324) and (hState = 351)) or
								((vState = 324) and (hState = 361)) or
								((vState = 324) and (hState = 366)) or
								((vState = 324) and (hState = 373)) or
								((vState = 324) and (hState = 384)) or
								((vState = 324) and (hState = 395)) or
								((vState = 324) and (hState = 401)) or
								((vState = 324) and (hState = 409)) or
								((vState = 324) and (hState = 418)) or
								((vState = 324) and (hState = 450)) or
								((vState = 324) and (hState = 481)) or
								((vState = 324) and (hState = 507)) or
								((vState = 324) and (hState = 519)) or
								((vState = 324) and (hState = 520)) or
								((vState = 324) and (hState = 521)) or
								((vState = 324) and (hState = 522)) or
								((vState = 324) and (hState = 528)) or
								((vState = 324) and (hState = 529)) or
								((vState = 324) and (hState = 530)) or
								((vState = 324) and (hState = 552)) or
								((vState = 324) and (hState = 576)) or
								((vState = 325) and (hState = 271)) or
								((vState = 325) and (hState = 292)) or
								((vState = 325) and (hState = 297)) or
								((vState = 325) and (hState = 304)) or
								((vState = 325) and (hState = 305)) or
								((vState = 325) and (hState = 319)) or
								((vState = 325) and (hState = 320)) or
								((vState = 325) and (hState = 361)) or
								((vState = 325) and (hState = 388)) or
								((vState = 325) and (hState = 395)) or
								((vState = 325) and (hState = 410)) or
								((vState = 325) and (hState = 519)) or
								((vState = 325) and (hState = 520)) or
								((vState = 325) and (hState = 528)) or
								((vState = 325) and (hState = 552)) or
								((vState = 326) and (hState = 271)) or
								((vState = 326) and (hState = 294)) or
								((vState = 326) and (hState = 295)) or
								((vState = 326) and (hState = 296)) or
								((vState = 326) and (hState = 297)) or
								((vState = 326) and (hState = 304)) or
								((vState = 326) and (hState = 305)) or
								((vState = 326) and (hState = 318)) or
								((vState = 326) and (hState = 319)) or
								((vState = 326) and (hState = 361)) or
								((vState = 326) and (hState = 386)) or
								((vState = 326) and (hState = 387)) or
								((vState = 326) and (hState = 388)) or
								((vState = 326) and (hState = 389)) or
								((vState = 326) and (hState = 394)) or
								((vState = 326) and (hState = 395)) or
								((vState = 326) and (hState = 411)) or
								((vState = 326) and (hState = 412)) or
								((vState = 326) and (hState = 413)) or
								((vState = 326) and (hState = 518)) or
								((vState = 326) and (hState = 541)) or
								((vState = 327) and (hState = 271)) or
								((vState = 327) and (hState = 294)) or
								((vState = 327) and (hState = 295)) or
								((vState = 327) and (hState = 296)) or
								((vState = 327) and (hState = 297)) or
								((vState = 327) and (hState = 304)) or
								((vState = 327) and (hState = 305)) or
								((vState = 327) and (hState = 318)) or
								((vState = 327) and (hState = 319)) or
								((vState = 327) and (hState = 339)) or
								((vState = 327) and (hState = 340)) or
								((vState = 327) and (hState = 361)) or
								((vState = 327) and (hState = 362)) or
								((vState = 327) and (hState = 386)) or
								((vState = 327) and (hState = 387)) or
								((vState = 327) and (hState = 388)) or
								((vState = 327) and (hState = 389)) or
								((vState = 327) and (hState = 390)) or
								((vState = 327) and (hState = 394)) or
								((vState = 327) and (hState = 395)) or
								((vState = 327) and (hState = 396)) or
								((vState = 327) and (hState = 411)) or
								((vState = 327) and (hState = 412)) or
								((vState = 327) and (hState = 413)) or
								((vState = 327) and (hState = 414)) or
								((vState = 327) and (hState = 415)) or
								((vState = 327) and (hState = 416)) or
								((vState = 327) and (hState = 422)) or
								((vState = 327) and (hState = 446)) or
								((vState = 327) and (hState = 453)) or
								((vState = 327) and (hState = 458)) or
								((vState = 327) and (hState = 512)) or
								((vState = 327) and (hState = 518)) or
								((vState = 327) and (hState = 527)) or
								((vState = 327) and (hState = 535)) or
								((vState = 327) and (hState = 541)) or
								((vState = 327) and (hState = 583)) or
								((vState = 327) and (hState = 584)) or
								((vState = 327) and (hState = 595)) or
								((vState = 327) and (hState = 596)) or
								((vState = 327) and (hState = 597)) or
								((vState = 328) and (hState = 294)) or
								((vState = 328) and (hState = 295)) or
								((vState = 328) and (hState = 296)) or
								((vState = 328) and (hState = 297)) or
								((vState = 328) and (hState = 298)) or
								((vState = 328) and (hState = 304)) or
								((vState = 328) and (hState = 317)) or
								((vState = 328) and (hState = 318)) or
								((vState = 328) and (hState = 319)) or
								((vState = 328) and (hState = 340)) or
								((vState = 328) and (hState = 361)) or
								((vState = 328) and (hState = 371)) or
								((vState = 328) and (hState = 388)) or
								((vState = 328) and (hState = 389)) or
								((vState = 328) and (hState = 390)) or
								((vState = 328) and (hState = 391)) or
								((vState = 328) and (hState = 392)) or
								((vState = 328) and (hState = 393)) or
								((vState = 328) and (hState = 394)) or
								((vState = 328) and (hState = 395)) or
								((vState = 328) and (hState = 412)) or
								((vState = 328) and (hState = 413)) or
								((vState = 328) and (hState = 417)) or
								((vState = 328) and (hState = 418)) or
								((vState = 328) and (hState = 422)) or
								((vState = 328) and (hState = 423)) or
								((vState = 328) and (hState = 424)) or
								((vState = 328) and (hState = 444)) or
								((vState = 328) and (hState = 445)) or
								((vState = 328) and (hState = 446)) or
								((vState = 328) and (hState = 454)) or
								((vState = 328) and (hState = 459)) or
								((vState = 328) and (hState = 475)) or
								((vState = 328) and (hState = 503)) or
								((vState = 328) and (hState = 511)) or
								((vState = 328) and (hState = 517)) or
								((vState = 328) and (hState = 537)) or
								((vState = 328) and (hState = 538)) or
								((vState = 328) and (hState = 539)) or
								((vState = 328) and (hState = 540)) or
								((vState = 328) and (hState = 541)) or
								((vState = 328) and (hState = 553)) or
								((vState = 328) and (hState = 587)) or
								((vState = 328) and (hState = 588)) or
								((vState = 328) and (hState = 589)) or
								((vState = 328) and (hState = 590)) or
								((vState = 328) and (hState = 591)) or
								((vState = 328) and (hState = 592)) or
								((vState = 328) and (hState = 593)) or
								((vState = 329) and (hState = 293)) or
								((vState = 329) and (hState = 297)) or
								((vState = 329) and (hState = 298)) or
								((vState = 329) and (hState = 299)) or
								((vState = 329) and (hState = 300)) or
								((vState = 329) and (hState = 304)) or
								((vState = 329) and (hState = 317)) or
								((vState = 329) and (hState = 318)) or
								((vState = 329) and (hState = 340)) or
								((vState = 329) and (hState = 341)) or
								((vState = 329) and (hState = 342)) or
								((vState = 329) and (hState = 347)) or
								((vState = 329) and (hState = 389)) or
								((vState = 329) and (hState = 390)) or
								((vState = 329) and (hState = 391)) or
								((vState = 329) and (hState = 392)) or
								((vState = 329) and (hState = 393)) or
								((vState = 329) and (hState = 412)) or
								((vState = 329) and (hState = 413)) or
								((vState = 329) and (hState = 421)) or
								((vState = 329) and (hState = 422)) or
								((vState = 329) and (hState = 423)) or
								((vState = 329) and (hState = 424)) or
								((vState = 329) and (hState = 425)) or
								((vState = 329) and (hState = 426)) or
								((vState = 329) and (hState = 427)) or
								((vState = 329) and (hState = 443)) or
								((vState = 329) and (hState = 455)) or
								((vState = 329) and (hState = 460)) or
								((vState = 329) and (hState = 497)) or
								((vState = 329) and (hState = 502)) or
								((vState = 329) and (hState = 525)) or
								((vState = 329) and (hState = 540)) or
								((vState = 329) and (hState = 541)) or
								((vState = 329) and (hState = 553)) or
								((vState = 330) and (hState = 297)) or
								((vState = 330) and (hState = 304)) or
								((vState = 330) and (hState = 340)) or
								((vState = 330) and (hState = 341)) or
								((vState = 330) and (hState = 389)) or
								((vState = 330) and (hState = 390)) or
								((vState = 330) and (hState = 391)) or
								((vState = 330) and (hState = 392)) or
								((vState = 330) and (hState = 412)) or
								((vState = 330) and (hState = 413)) or
								((vState = 330) and (hState = 423)) or
								((vState = 330) and (hState = 424)) or
								((vState = 330) and (hState = 425)) or
								((vState = 330) and (hState = 426)) or
								((vState = 330) and (hState = 427)) or
								((vState = 330) and (hState = 525)) or
								((vState = 330) and (hState = 553)) or
								((vState = 331) and (hState = 297)) or
								((vState = 331) and (hState = 303)) or
								((vState = 331) and (hState = 304)) or
								((vState = 331) and (hState = 315)) or
								((vState = 331) and (hState = 340)) or
								((vState = 331) and (hState = 341)) or
								((vState = 331) and (hState = 359)) or
								((vState = 331) and (hState = 389)) or
								((vState = 331) and (hState = 390)) or
								((vState = 331) and (hState = 391)) or
								((vState = 331) and (hState = 392)) or
								((vState = 331) and (hState = 393)) or
								((vState = 331) and (hState = 412)) or
								((vState = 331) and (hState = 413)) or
								((vState = 331) and (hState = 427)) or
								((vState = 331) and (hState = 428)) or
								((vState = 331) and (hState = 429)) or
								((vState = 331) and (hState = 513)) or
								((vState = 331) and (hState = 553)) or
								((vState = 332) and (hState = 297)) or
								((vState = 332) and (hState = 303)) or
								((vState = 332) and (hState = 304)) or
								((vState = 332) and (hState = 305)) or
								((vState = 332) and (hState = 315)) or
								((vState = 332) and (hState = 340)) or
								((vState = 332) and (hState = 341)) or
								((vState = 332) and (hState = 346)) or
								((vState = 332) and (hState = 356)) or
								((vState = 332) and (hState = 368)) or
								((vState = 332) and (hState = 389)) or
								((vState = 332) and (hState = 390)) or
								((vState = 332) and (hState = 391)) or
								((vState = 332) and (hState = 392)) or
								((vState = 332) and (hState = 393)) or
								((vState = 332) and (hState = 394)) or
								((vState = 332) and (hState = 412)) or
								((vState = 332) and (hState = 413)) or
								((vState = 332) and (hState = 427)) or
								((vState = 332) and (hState = 428)) or
								((vState = 332) and (hState = 429)) or
								((vState = 332) and (hState = 430)) or
								((vState = 332) and (hState = 431)) or
								((vState = 332) and (hState = 432)) or
								((vState = 332) and (hState = 458)) or
								((vState = 332) and (hState = 469)) or
								((vState = 332) and (hState = 507)) or
								((vState = 332) and (hState = 512)) or
								((vState = 332) and (hState = 513)) or
								((vState = 332) and (hState = 527)) or
								((vState = 332) and (hState = 528)) or
								((vState = 332) and (hState = 553)) or
								((vState = 333) and (hState = 290)) or
								((vState = 333) and (hState = 297)) or
								((vState = 333) and (hState = 303)) or
								((vState = 333) and (hState = 304)) or
								((vState = 333) and (hState = 305)) or
								((vState = 333) and (hState = 306)) or
								((vState = 333) and (hState = 307)) or
								((vState = 333) and (hState = 308)) or
								((vState = 333) and (hState = 314)) or
								((vState = 333) and (hState = 315)) or
								((vState = 333) and (hState = 340)) or
								((vState = 333) and (hState = 345)) or
								((vState = 333) and (hState = 355)) or
								((vState = 333) and (hState = 386)) or
								((vState = 333) and (hState = 387)) or
								((vState = 333) and (hState = 391)) or
								((vState = 333) and (hState = 392)) or
								((vState = 333) and (hState = 393)) or
								((vState = 333) and (hState = 394)) or
								((vState = 333) and (hState = 395)) or
								((vState = 333) and (hState = 412)) or
								((vState = 333) and (hState = 413)) or
								((vState = 333) and (hState = 414)) or
								((vState = 333) and (hState = 429)) or
								((vState = 333) and (hState = 430)) or
								((vState = 333) and (hState = 431)) or
								((vState = 333) and (hState = 432)) or
								((vState = 333) and (hState = 433)) or
								((vState = 333) and (hState = 434)) or
								((vState = 333) and (hState = 439)) or
								((vState = 333) and (hState = 459)) or
								((vState = 333) and (hState = 466)) or
								((vState = 333) and (hState = 467)) or
								((vState = 333) and (hState = 506)) or
								((vState = 333) and (hState = 512)) or
								((vState = 333) and (hState = 523)) or
								((vState = 333) and (hState = 529)) or
								((vState = 333) and (hState = 530)) or
								((vState = 333) and (hState = 565)) or
								((vState = 334) and (hState = 289)) or
								((vState = 334) and (hState = 309)) or
								((vState = 334) and (hState = 310)) or
								((vState = 334) and (hState = 311)) or
								((vState = 334) and (hState = 312)) or
								((vState = 334) and (hState = 313)) or
								((vState = 334) and (hState = 314)) or
								((vState = 334) and (hState = 340)) or
								((vState = 334) and (hState = 367)) or
								((vState = 334) and (hState = 384)) or
								((vState = 334) and (hState = 391)) or
								((vState = 334) and (hState = 392)) or
								((vState = 334) and (hState = 393)) or
								((vState = 334) and (hState = 394)) or
								((vState = 334) and (hState = 395)) or
								((vState = 334) and (hState = 396)) or
								((vState = 334) and (hState = 412)) or
								((vState = 334) and (hState = 416)) or
								((vState = 334) and (hState = 433)) or
								((vState = 334) and (hState = 434)) or
								((vState = 334) and (hState = 435)) or
								((vState = 334) and (hState = 436)) or
								((vState = 334) and (hState = 437)) or
								((vState = 334) and (hState = 438)) or
								((vState = 334) and (hState = 439)) or
								((vState = 334) and (hState = 460)) or
								((vState = 334) and (hState = 464)) or
								((vState = 334) and (hState = 465)) or
								((vState = 334) and (hState = 501)) or
								((vState = 334) and (hState = 511)) or
								((vState = 334) and (hState = 522)) or
								((vState = 334) and (hState = 530)) or
								((vState = 334) and (hState = 531)) or
								((vState = 334) and (hState = 532)) or
								((vState = 334) and (hState = 552)) or
								((vState = 334) and (hState = 562)) or
								((vState = 334) and (hState = 563)) or
								((vState = 334) and (hState = 564)) or
								((vState = 334) and (hState = 565)) or
								((vState = 335) and (hState = 312)) or
								((vState = 335) and (hState = 313)) or
								((vState = 335) and (hState = 314)) or
								((vState = 335) and (hState = 340)) or
								((vState = 335) and (hState = 395)) or
								((vState = 335) and (hState = 396)) or
								((vState = 335) and (hState = 412)) or
								((vState = 335) and (hState = 436)) or
								((vState = 335) and (hState = 437)) or
								((vState = 335) and (hState = 438)) or
								((vState = 335) and (hState = 439)) or
								((vState = 335) and (hState = 464)) or
								((vState = 335) and (hState = 465)) or
								((vState = 335) and (hState = 511)) or
								((vState = 335) and (hState = 532)) or
								((vState = 335) and (hState = 533)) or
								((vState = 336) and (hState = 312)) or
								((vState = 336) and (hState = 313)) or
								((vState = 336) and (hState = 314)) or
								((vState = 336) and (hState = 366)) or
								((vState = 336) and (hState = 396)) or
								((vState = 336) and (hState = 397)) or
								((vState = 336) and (hState = 398)) or
								((vState = 336) and (hState = 436)) or
								((vState = 336) and (hState = 437)) or
								((vState = 336) and (hState = 438)) or
								((vState = 336) and (hState = 439)) or
								((vState = 336) and (hState = 502)) or
								((vState = 336) and (hState = 503)) or
								((vState = 336) and (hState = 534)) or
								((vState = 336) and (hState = 535)) or
								((vState = 336) and (hState = 551)) or
								((vState = 337) and (hState = 287)) or
								((vState = 337) and (hState = 312)) or
								((vState = 337) and (hState = 365)) or
								((vState = 337) and (hState = 390)) or
								((vState = 337) and (hState = 397)) or
								((vState = 337) and (hState = 398)) or
								((vState = 337) and (hState = 441)) or
								((vState = 337) and (hState = 442)) or
								((vState = 337) and (hState = 443)) or
								((vState = 337) and (hState = 502)) or
								((vState = 337) and (hState = 503)) or
								((vState = 337) and (hState = 535)) or
								((vState = 337) and (hState = 536)) or
								((vState = 337) and (hState = 537)) or
								((vState = 337) and (hState = 538)) or
								((vState = 337) and (hState = 539)) or
								((vState = 337) and (hState = 551)) or
								((vState = 337) and (hState = 557)) or
								((vState = 338) and (hState = 317)) or
								((vState = 338) and (hState = 318)) or
								((vState = 338) and (hState = 360)) or
								((vState = 338) and (hState = 361)) or
								((vState = 338) and (hState = 362)) or
								((vState = 338) and (hState = 363)) or
								((vState = 338) and (hState = 364)) or
								((vState = 338) and (hState = 378)) or
								((vState = 338) and (hState = 390)) or
								((vState = 338) and (hState = 397)) or
								((vState = 338) and (hState = 398)) or
								((vState = 338) and (hState = 411)) or
								((vState = 338) and (hState = 418)) or
								((vState = 338) and (hState = 434)) or
								((vState = 338) and (hState = 442)) or
								((vState = 338) and (hState = 443)) or
								((vState = 338) and (hState = 444)) or
								((vState = 338) and (hState = 445)) or
								((vState = 338) and (hState = 446)) or
								((vState = 338) and (hState = 490)) or
								((vState = 338) and (hState = 502)) or
								((vState = 338) and (hState = 503)) or
								((vState = 338) and (hState = 504)) or
								((vState = 338) and (hState = 508)) or
								((vState = 338) and (hState = 519)) or
								((vState = 338) and (hState = 536)) or
								((vState = 338) and (hState = 537)) or
								((vState = 338) and (hState = 538)) or
								((vState = 338) and (hState = 539)) or
								((vState = 338) and (hState = 540)) or
								((vState = 338) and (hState = 541)) or
								((vState = 338) and (hState = 550)) or
								((vState = 338) and (hState = 551)) or
								((vState = 338) and (hState = 555)) or
								((vState = 338) and (hState = 556)) or
								((vState = 339) and (hState = 267)) or
								((vState = 339) and (hState = 310)) or
								((vState = 339) and (hState = 319)) or
								((vState = 339) and (hState = 320)) or
								((vState = 339) and (hState = 338)) or
								((vState = 339) and (hState = 339)) or
								((vState = 339) and (hState = 340)) or
								((vState = 339) and (hState = 341)) or
								((vState = 339) and (hState = 347)) or
								((vState = 339) and (hState = 348)) or
								((vState = 339) and (hState = 355)) or
								((vState = 339) and (hState = 356)) or
								((vState = 339) and (hState = 357)) or
								((vState = 339) and (hState = 358)) or
								((vState = 339) and (hState = 359)) or
								((vState = 339) and (hState = 360)) or
								((vState = 339) and (hState = 361)) or
								((vState = 339) and (hState = 362)) or
								((vState = 339) and (hState = 363)) or
								((vState = 339) and (hState = 378)) or
								((vState = 339) and (hState = 397)) or
								((vState = 339) and (hState = 398)) or
								((vState = 339) and (hState = 399)) or
								((vState = 339) and (hState = 400)) or
								((vState = 339) and (hState = 411)) or
								((vState = 339) and (hState = 433)) or
								((vState = 339) and (hState = 443)) or
								((vState = 339) and (hState = 447)) or
								((vState = 339) and (hState = 448)) or
								((vState = 339) and (hState = 501)) or
								((vState = 339) and (hState = 506)) or
								((vState = 339) and (hState = 507)) or
								((vState = 339) and (hState = 508)) or
								((vState = 339) and (hState = 518)) or
								((vState = 339) and (hState = 537)) or
								((vState = 339) and (hState = 538)) or
								((vState = 339) and (hState = 539)) or
								((vState = 339) and (hState = 540)) or
								((vState = 339) and (hState = 541)) or
								((vState = 339) and (hState = 542)) or
								((vState = 339) and (hState = 543)) or
								((vState = 339) and (hState = 550)) or
								((vState = 339) and (hState = 551)) or
								((vState = 339) and (hState = 552)) or
								((vState = 339) and (hState = 553)) or
								((vState = 340) and (hState = 267)) or
								((vState = 340) and (hState = 295)) or
								((vState = 340) and (hState = 310)) or
								((vState = 340) and (hState = 338)) or
								((vState = 340) and (hState = 339)) or
								((vState = 340) and (hState = 340)) or
								((vState = 340) and (hState = 347)) or
								((vState = 340) and (hState = 348)) or
								((vState = 340) and (hState = 349)) or
								((vState = 340) and (hState = 360)) or
								((vState = 340) and (hState = 361)) or
								((vState = 340) and (hState = 362)) or
								((vState = 340) and (hState = 363)) or
								((vState = 340) and (hState = 378)) or
								((vState = 340) and (hState = 397)) or
								((vState = 340) and (hState = 411)) or
								((vState = 340) and (hState = 443)) or
								((vState = 340) and (hState = 506)) or
								((vState = 340) and (hState = 507)) or
								((vState = 340) and (hState = 508)) or
								((vState = 340) and (hState = 540)) or
								((vState = 340) and (hState = 541)) or
								((vState = 340) and (hState = 542)) or
								((vState = 340) and (hState = 550)) or
								((vState = 340) and (hState = 551)) or
								((vState = 341) and (hState = 267)) or
								((vState = 341) and (hState = 294)) or
								((vState = 341) and (hState = 295)) or
								((vState = 341) and (hState = 337)) or
								((vState = 341) and (hState = 338)) or
								((vState = 341) and (hState = 339)) or
								((vState = 341) and (hState = 340)) or
								((vState = 341) and (hState = 346)) or
								((vState = 341) and (hState = 347)) or
								((vState = 341) and (hState = 360)) or
								((vState = 341) and (hState = 361)) or
								((vState = 341) and (hState = 362)) or
								((vState = 341) and (hState = 378)) or
								((vState = 341) and (hState = 389)) or
								((vState = 341) and (hState = 411)) or
								((vState = 341) and (hState = 443)) or
								((vState = 341) and (hState = 506)) or
								((vState = 341) and (hState = 507)) or
								((vState = 341) and (hState = 508)) or
								((vState = 341) and (hState = 540)) or
								((vState = 341) and (hState = 541)) or
								((vState = 341) and (hState = 542)) or
								((vState = 341) and (hState = 546)) or
								((vState = 341) and (hState = 547)) or
								((vState = 341) and (hState = 548)) or
								((vState = 341) and (hState = 549)) or
								((vState = 341) and (hState = 550)) or
								((vState = 341) and (hState = 551)) or
								((vState = 342) and (hState = 294)) or
								((vState = 342) and (hState = 295)) or
								((vState = 342) and (hState = 299)) or
								((vState = 342) and (hState = 307)) or
								((vState = 342) and (hState = 308)) or
								((vState = 342) and (hState = 309)) or
								((vState = 342) and (hState = 324)) or
								((vState = 342) and (hState = 336)) or
								((vState = 342) and (hState = 337)) or
								((vState = 342) and (hState = 338)) or
								((vState = 342) and (hState = 339)) or
								((vState = 342) and (hState = 340)) or
								((vState = 342) and (hState = 360)) or
								((vState = 342) and (hState = 361)) or
								((vState = 342) and (hState = 506)) or
								((vState = 342) and (hState = 540)) or
								((vState = 342) and (hState = 541)) or
								((vState = 342) and (hState = 542)) or
								((vState = 342) and (hState = 546)) or
								((vState = 342) and (hState = 547)) or
								((vState = 342) and (hState = 548)) or
								((vState = 342) and (hState = 549)) or
								((vState = 342) and (hState = 550)) or
								((vState = 342) and (hState = 551)) or
								((vState = 343) and (hState = 266)) or
								((vState = 343) and (hState = 282)) or
								((vState = 343) and (hState = 294)) or
								((vState = 343) and (hState = 295)) or
								((vState = 343) and (hState = 296)) or
								((vState = 343) and (hState = 297)) or
								((vState = 343) and (hState = 298)) or
								((vState = 343) and (hState = 299)) or
								((vState = 343) and (hState = 307)) or
								((vState = 343) and (hState = 308)) or
								((vState = 343) and (hState = 309)) or
								((vState = 343) and (hState = 324)) or
								((vState = 343) and (hState = 336)) or
								((vState = 343) and (hState = 337)) or
								((vState = 343) and (hState = 338)) or
								((vState = 343) and (hState = 339)) or
								((vState = 343) and (hState = 340)) or
								((vState = 343) and (hState = 341)) or
								((vState = 343) and (hState = 342)) or
								((vState = 343) and (hState = 360)) or
								((vState = 343) and (hState = 361)) or
								((vState = 343) and (hState = 429)) or
								((vState = 343) and (hState = 455)) or
								((vState = 343) and (hState = 471)) or
								((vState = 343) and (hState = 485)) or
								((vState = 343) and (hState = 497)) or
								((vState = 343) and (hState = 505)) or
								((vState = 343) and (hState = 506)) or
								((vState = 343) and (hState = 511)) or
								((vState = 343) and (hState = 536)) or
								((vState = 343) and (hState = 537)) or
								((vState = 343) and (hState = 538)) or
								((vState = 343) and (hState = 539)) or
								((vState = 343) and (hState = 540)) or
								((vState = 343) and (hState = 541)) or
								((vState = 343) and (hState = 542)) or
								((vState = 343) and (hState = 543)) or
								((vState = 343) and (hState = 544)) or
								((vState = 343) and (hState = 545)) or
								((vState = 343) and (hState = 546)) or
								((vState = 343) and (hState = 547)) or
								((vState = 343) and (hState = 548)) or
								((vState = 343) and (hState = 549)) or
								((vState = 343) and (hState = 550)) or
								((vState = 343) and (hState = 551)) or
								((vState = 343) and (hState = 573)) or
								((vState = 343) and (hState = 574)) or
								((vState = 343) and (hState = 575)) or
								((vState = 343) and (hState = 576)) or
								((vState = 343) and (hState = 577)) or
								((vState = 343) and (hState = 581)) or
								((vState = 343) and (hState = 582)) or
								((vState = 343) and (hState = 583)) or
								((vState = 343) and (hState = 584)) or
								((vState = 343) and (hState = 585)) or
								((vState = 343) and (hState = 586)) or
								((vState = 343) and (hState = 587)) or
								((vState = 343) and (hState = 588)) or
								((vState = 343) and (hState = 589)) or
								((vState = 343) and (hState = 590)) or
								((vState = 344) and (hState = 266)) or
								((vState = 344) and (hState = 281)) or
								((vState = 344) and (hState = 294)) or
								((vState = 344) and (hState = 295)) or
								((vState = 344) and (hState = 296)) or
								((vState = 344) and (hState = 297)) or
								((vState = 344) and (hState = 298)) or
								((vState = 344) and (hState = 299)) or
								((vState = 344) and (hState = 307)) or
								((vState = 344) and (hState = 308)) or
								((vState = 344) and (hState = 309)) or
								((vState = 344) and (hState = 310)) or
								((vState = 344) and (hState = 311)) or
								((vState = 344) and (hState = 312)) or
								((vState = 344) and (hState = 313)) or
								((vState = 344) and (hState = 314)) or
								((vState = 344) and (hState = 315)) or
								((vState = 344) and (hState = 316)) or
								((vState = 344) and (hState = 317)) or
								((vState = 344) and (hState = 318)) or
								((vState = 344) and (hState = 324)) or
								((vState = 344) and (hState = 335)) or
								((vState = 344) and (hState = 339)) or
								((vState = 344) and (hState = 340)) or
								((vState = 344) and (hState = 341)) or
								((vState = 344) and (hState = 360)) or
								((vState = 344) and (hState = 361)) or
								((vState = 344) and (hState = 379)) or
								((vState = 344) and (hState = 388)) or
								((vState = 344) and (hState = 422)) or
								((vState = 344) and (hState = 428)) or
								((vState = 344) and (hState = 429)) or
								((vState = 344) and (hState = 448)) or
								((vState = 344) and (hState = 458)) or
								((vState = 344) and (hState = 459)) or
								((vState = 344) and (hState = 496)) or
								((vState = 344) and (hState = 497)) or
								((vState = 344) and (hState = 503)) or
								((vState = 344) and (hState = 504)) or
								((vState = 344) and (hState = 505)) or
								((vState = 344) and (hState = 506)) or
								((vState = 344) and (hState = 512)) or
								((vState = 344) and (hState = 513)) or
								((vState = 344) and (hState = 514)) or
								((vState = 344) and (hState = 534)) or
								((vState = 344) and (hState = 540)) or
								((vState = 344) and (hState = 541)) or
								((vState = 344) and (hState = 542)) or
								((vState = 344) and (hState = 543)) or
								((vState = 344) and (hState = 544)) or
								((vState = 344) and (hState = 545)) or
								((vState = 344) and (hState = 546)) or
								((vState = 344) and (hState = 547)) or
								((vState = 344) and (hState = 552)) or
								((vState = 344) and (hState = 553)) or
								((vState = 344) and (hState = 554)) or
								((vState = 344) and (hState = 555)) or
								((vState = 344) and (hState = 556)) or
								((vState = 344) and (hState = 557)) or
								((vState = 344) and (hState = 558)) or
								((vState = 344) and (hState = 559)) or
								((vState = 344) and (hState = 560)) or
								((vState = 344) and (hState = 561)) or
								((vState = 344) and (hState = 562)) or
								((vState = 344) and (hState = 563)) or
								((vState = 344) and (hState = 564)) or
								((vState = 344) and (hState = 565)) or
								((vState = 344) and (hState = 566)) or
								((vState = 344) and (hState = 567)) or
								((vState = 344) and (hState = 568)) or
								((vState = 344) and (hState = 569)) or
								((vState = 345) and (hState = 266)) or
								((vState = 345) and (hState = 294)) or
								((vState = 345) and (hState = 295)) or
								((vState = 345) and (hState = 296)) or
								((vState = 345) and (hState = 297)) or
								((vState = 345) and (hState = 298)) or
								((vState = 345) and (hState = 299)) or
								((vState = 345) and (hState = 300)) or
								((vState = 345) and (hState = 320)) or
								((vState = 345) and (hState = 321)) or
								((vState = 345) and (hState = 322)) or
								((vState = 345) and (hState = 323)) or
								((vState = 345) and (hState = 324)) or
								((vState = 345) and (hState = 325)) or
								((vState = 345) and (hState = 326)) or
								((vState = 345) and (hState = 327)) or
								((vState = 345) and (hState = 335)) or
								((vState = 345) and (hState = 339)) or
								((vState = 345) and (hState = 340)) or
								((vState = 345) and (hState = 379)) or
								((vState = 345) and (hState = 388)) or
								((vState = 345) and (hState = 423)) or
								((vState = 345) and (hState = 424)) or
								((vState = 345) and (hState = 425)) or
								((vState = 345) and (hState = 426)) or
								((vState = 345) and (hState = 427)) or
								((vState = 345) and (hState = 428)) or
								((vState = 345) and (hState = 429)) or
								((vState = 345) and (hState = 448)) or
								((vState = 345) and (hState = 460)) or
								((vState = 345) and (hState = 461)) or
								((vState = 345) and (hState = 474)) or
								((vState = 345) and (hState = 490)) or
								((vState = 345) and (hState = 491)) or
								((vState = 345) and (hState = 492)) or
								((vState = 345) and (hState = 493)) or
								((vState = 345) and (hState = 494)) or
								((vState = 345) and (hState = 495)) or
								((vState = 345) and (hState = 496)) or
								((vState = 345) and (hState = 497)) or
								((vState = 345) and (hState = 498)) or
								((vState = 345) and (hState = 499)) or
								((vState = 345) and (hState = 500)) or
								((vState = 345) and (hState = 501)) or
								((vState = 345) and (hState = 502)) or
								((vState = 345) and (hState = 503)) or
								((vState = 345) and (hState = 504)) or
								((vState = 345) and (hState = 513)) or
								((vState = 345) and (hState = 514)) or
								((vState = 345) and (hState = 530)) or
								((vState = 345) and (hState = 531)) or
								((vState = 345) and (hState = 540)) or
								((vState = 345) and (hState = 541)) or
								((vState = 345) and (hState = 545)) or
								((vState = 345) and (hState = 546)) or
								((vState = 345) and (hState = 547)) or
								((vState = 345) and (hState = 553)) or
								((vState = 345) and (hState = 554)) or
								((vState = 345) and (hState = 555)) or
								((vState = 345) and (hState = 556)) or
								((vState = 345) and (hState = 557)) or
								((vState = 345) and (hState = 558)) or
								((vState = 345) and (hState = 559)) or
								((vState = 346) and (hState = 294)) or
								((vState = 346) and (hState = 295)) or
								((vState = 346) and (hState = 296)) or
								((vState = 346) and (hState = 297)) or
								((vState = 346) and (hState = 298)) or
								((vState = 346) and (hState = 325)) or
								((vState = 346) and (hState = 326)) or
								((vState = 346) and (hState = 335)) or
								((vState = 346) and (hState = 339)) or
								((vState = 346) and (hState = 340)) or
								((vState = 346) and (hState = 425)) or
								((vState = 346) and (hState = 426)) or
								((vState = 346) and (hState = 427)) or
								((vState = 346) and (hState = 428)) or
								((vState = 346) and (hState = 429)) or
								((vState = 346) and (hState = 448)) or
								((vState = 346) and (hState = 460)) or
								((vState = 346) and (hState = 461)) or
								((vState = 346) and (hState = 474)) or
								((vState = 346) and (hState = 490)) or
								((vState = 346) and (hState = 491)) or
								((vState = 346) and (hState = 492)) or
								((vState = 346) and (hState = 493)) or
								((vState = 346) and (hState = 503)) or
								((vState = 346) and (hState = 504)) or
								((vState = 346) and (hState = 513)) or
								((vState = 346) and (hState = 514)) or
								((vState = 346) and (hState = 545)) or
								((vState = 346) and (hState = 556)) or
								((vState = 346) and (hState = 557)) or
								((vState = 346) and (hState = 558)) or
								((vState = 346) and (hState = 559)) or
								((vState = 347) and (hState = 294)) or
								((vState = 347) and (hState = 295)) or
								((vState = 347) and (hState = 296)) or
								((vState = 347) and (hState = 297)) or
								((vState = 347) and (hState = 298)) or
								((vState = 347) and (hState = 303)) or
								((vState = 347) and (hState = 304)) or
								((vState = 347) and (hState = 305)) or
								((vState = 347) and (hState = 306)) or
								((vState = 347) and (hState = 326)) or
								((vState = 347) and (hState = 334)) or
								((vState = 347) and (hState = 335)) or
								((vState = 347) and (hState = 336)) or
								((vState = 347) and (hState = 337)) or
								((vState = 347) and (hState = 407)) or
								((vState = 347) and (hState = 448)) or
								((vState = 347) and (hState = 460)) or
								((vState = 347) and (hState = 461)) or
								((vState = 347) and (hState = 462)) or
								((vState = 347) and (hState = 463)) or
								((vState = 347) and (hState = 464)) or
								((vState = 347) and (hState = 476)) or
								((vState = 347) and (hState = 480)) or
								((vState = 347) and (hState = 481)) or
								((vState = 347) and (hState = 490)) or
								((vState = 347) and (hState = 491)) or
								((vState = 347) and (hState = 492)) or
								((vState = 347) and (hState = 493)) or
								((vState = 347) and (hState = 503)) or
								((vState = 347) and (hState = 557)) or
								((vState = 347) and (hState = 558)) or
								((vState = 348) and (hState = 294)) or
								((vState = 348) and (hState = 295)) or
								((vState = 348) and (hState = 296)) or
								((vState = 348) and (hState = 297)) or
								((vState = 348) and (hState = 298)) or
								((vState = 348) and (hState = 303)) or
								((vState = 348) and (hState = 304)) or
								((vState = 348) and (hState = 305)) or
								((vState = 348) and (hState = 306)) or
								((vState = 348) and (hState = 326)) or
								((vState = 348) and (hState = 334)) or
								((vState = 348) and (hState = 335)) or
								((vState = 348) and (hState = 336)) or
								((vState = 348) and (hState = 337)) or
								((vState = 348) and (hState = 341)) or
								((vState = 348) and (hState = 342)) or
								((vState = 348) and (hState = 343)) or
								((vState = 348) and (hState = 344)) or
								((vState = 348) and (hState = 345)) or
								((vState = 348) and (hState = 346)) or
								((vState = 348) and (hState = 347)) or
								((vState = 348) and (hState = 348)) or
								((vState = 348) and (hState = 358)) or
								((vState = 348) and (hState = 386)) or
								((vState = 348) and (hState = 387)) or
								((vState = 348) and (hState = 407)) or
								((vState = 348) and (hState = 431)) or
								((vState = 348) and (hState = 432)) or
								((vState = 348) and (hState = 433)) or
								((vState = 348) and (hState = 448)) or
								((vState = 348) and (hState = 459)) or
								((vState = 348) and (hState = 460)) or
								((vState = 348) and (hState = 461)) or
								((vState = 348) and (hState = 462)) or
								((vState = 348) and (hState = 463)) or
								((vState = 348) and (hState = 464)) or
								((vState = 348) and (hState = 465)) or
								((vState = 348) and (hState = 466)) or
								((vState = 348) and (hState = 467)) or
								((vState = 348) and (hState = 468)) or
								((vState = 348) and (hState = 469)) or
								((vState = 348) and (hState = 470)) or
								((vState = 348) and (hState = 471)) or
								((vState = 348) and (hState = 476)) or
								((vState = 348) and (hState = 480)) or
								((vState = 348) and (hState = 481)) or
								((vState = 348) and (hState = 490)) or
								((vState = 348) and (hState = 491)) or
								((vState = 348) and (hState = 492)) or
								((vState = 348) and (hState = 493)) or
								((vState = 348) and (hState = 503)) or
								((vState = 348) and (hState = 512)) or
								((vState = 348) and (hState = 525)) or
								((vState = 348) and (hState = 535)) or
								((vState = 348) and (hState = 536)) or
								((vState = 348) and (hState = 551)) or
								((vState = 348) and (hState = 557)) or
								((vState = 348) and (hState = 558)) or
								((vState = 348) and (hState = 562)) or
								((vState = 348) and (hState = 563)) or
								((vState = 348) and (hState = 564)) or
								((vState = 349) and (hState = 294)) or
								((vState = 349) and (hState = 295)) or
								((vState = 349) and (hState = 296)) or
								((vState = 349) and (hState = 297)) or
								((vState = 349) and (hState = 298)) or
								((vState = 349) and (hState = 303)) or
								((vState = 349) and (hState = 326)) or
								((vState = 349) and (hState = 334)) or
								((vState = 349) and (hState = 335)) or
								((vState = 349) and (hState = 336)) or
								((vState = 349) and (hState = 337)) or
								((vState = 349) and (hState = 351)) or
								((vState = 349) and (hState = 352)) or
								((vState = 349) and (hState = 353)) or
								((vState = 349) and (hState = 354)) or
								((vState = 349) and (hState = 355)) or
								((vState = 349) and (hState = 356)) or
								((vState = 349) and (hState = 357)) or
								((vState = 349) and (hState = 358)) or
								((vState = 349) and (hState = 386)) or
								((vState = 349) and (hState = 387)) or
								((vState = 349) and (hState = 400)) or
								((vState = 349) and (hState = 407)) or
								((vState = 349) and (hState = 408)) or
								((vState = 349) and (hState = 423)) or
								((vState = 349) and (hState = 436)) or
								((vState = 349) and (hState = 437)) or
								((vState = 349) and (hState = 448)) or
								((vState = 349) and (hState = 469)) or
								((vState = 349) and (hState = 470)) or
								((vState = 349) and (hState = 471)) or
								((vState = 349) and (hState = 476)) or
								((vState = 349) and (hState = 480)) or
								((vState = 349) and (hState = 490)) or
								((vState = 349) and (hState = 491)) or
								((vState = 349) and (hState = 492)) or
								((vState = 349) and (hState = 493)) or
								((vState = 349) and (hState = 511)) or
								((vState = 349) and (hState = 517)) or
								((vState = 349) and (hState = 522)) or
								((vState = 349) and (hState = 523)) or
								((vState = 349) and (hState = 532)) or
								((vState = 349) and (hState = 533)) or
								((vState = 349) and (hState = 534)) or
								((vState = 349) and (hState = 553)) or
								((vState = 349) and (hState = 557)) or
								((vState = 349) and (hState = 558)) or
								((vState = 349) and (hState = 563)) or
								((vState = 349) and (hState = 564)) or
								((vState = 349) and (hState = 565)) or
								((vState = 349) and (hState = 566)) or
								((vState = 349) and (hState = 567)) or
								((vState = 350) and (hState = 294)) or
								((vState = 350) and (hState = 295)) or
								((vState = 350) and (hState = 299)) or
								((vState = 350) and (hState = 308)) or
								((vState = 350) and (hState = 333)) or
								((vState = 350) and (hState = 334)) or
								((vState = 350) and (hState = 356)) or
								((vState = 350) and (hState = 357)) or
								((vState = 350) and (hState = 358)) or
								((vState = 350) and (hState = 359)) or
								((vState = 350) and (hState = 360)) or
								((vState = 350) and (hState = 361)) or
								((vState = 350) and (hState = 362)) or
								((vState = 350) and (hState = 363)) or
								((vState = 350) and (hState = 364)) or
								((vState = 350) and (hState = 365)) or
								((vState = 350) and (hState = 366)) or
								((vState = 350) and (hState = 367)) or
								((vState = 350) and (hState = 368)) or
								((vState = 350) and (hState = 369)) or
								((vState = 350) and (hState = 400)) or
								((vState = 350) and (hState = 406)) or
								((vState = 350) and (hState = 422)) or
								((vState = 350) and (hState = 439)) or
								((vState = 350) and (hState = 440)) or
								((vState = 350) and (hState = 448)) or
								((vState = 350) and (hState = 471)) or
								((vState = 350) and (hState = 476)) or
								((vState = 350) and (hState = 477)) or
								((vState = 350) and (hState = 478)) or
								((vState = 350) and (hState = 489)) or
								((vState = 350) and (hState = 490)) or
								((vState = 350) and (hState = 491)) or
								((vState = 350) and (hState = 496)) or
								((vState = 350) and (hState = 502)) or
								((vState = 350) and (hState = 517)) or
								((vState = 350) and (hState = 518)) or
								((vState = 350) and (hState = 519)) or
								((vState = 350) and (hState = 520)) or
								((vState = 350) and (hState = 530)) or
								((vState = 350) and (hState = 531)) or
								((vState = 350) and (hState = 542)) or
								((vState = 350) and (hState = 555)) or
								((vState = 350) and (hState = 556)) or
								((vState = 350) and (hState = 557)) or
								((vState = 350) and (hState = 558)) or
								((vState = 350) and (hState = 559)) or
								((vState = 350) and (hState = 563)) or
								((vState = 350) and (hState = 567)) or
								((vState = 350) and (hState = 568)) or
								((vState = 350) and (hState = 569)) or
								((vState = 351) and (hState = 294)) or
								((vState = 351) and (hState = 295)) or
								((vState = 351) and (hState = 308)) or
								((vState = 351) and (hState = 357)) or
								((vState = 351) and (hState = 358)) or
								((vState = 351) and (hState = 439)) or
								((vState = 351) and (hState = 448)) or
								((vState = 351) and (hState = 476)) or
								((vState = 351) and (hState = 477)) or
								((vState = 351) and (hState = 489)) or
								((vState = 351) and (hState = 490)) or
								((vState = 351) and (hState = 517)) or
								((vState = 351) and (hState = 518)) or
								((vState = 351) and (hState = 519)) or
								((vState = 351) and (hState = 520)) or
								((vState = 351) and (hState = 557)) or
								((vState = 351) and (hState = 558)) or
								((vState = 351) and (hState = 559)) or
								((vState = 351) and (hState = 560)) or
								((vState = 351) and (hState = 563)) or
								((vState = 351) and (hState = 569)) or
								((vState = 352) and (hState = 294)) or
								((vState = 352) and (hState = 295)) or
								((vState = 352) and (hState = 301)) or
								((vState = 352) and (hState = 308)) or
								((vState = 352) and (hState = 331)) or
								((vState = 352) and (hState = 358)) or
								((vState = 352) and (hState = 382)) or
								((vState = 352) and (hState = 385)) or
								((vState = 352) and (hState = 439)) or
								((vState = 352) and (hState = 448)) or
								((vState = 352) and (hState = 476)) or
								((vState = 352) and (hState = 477)) or
								((vState = 352) and (hState = 520)) or
								((vState = 352) and (hState = 558)) or
								((vState = 352) and (hState = 559)) or
								((vState = 352) and (hState = 560)) or
								((vState = 352) and (hState = 561)) or
								((vState = 352) and (hState = 562)) or
								((vState = 352) and (hState = 563)) or
								((vState = 352) and (hState = 572)) or
								((vState = 352) and (hState = 573)) or
								((vState = 353) and (hState = 293)) or
								((vState = 353) and (hState = 294)) or
								((vState = 353) and (hState = 295)) or
								((vState = 353) and (hState = 301)) or
								((vState = 353) and (hState = 308)) or
								((vState = 353) and (hState = 328)) or
								((vState = 353) and (hState = 329)) or
								((vState = 353) and (hState = 330)) or
								((vState = 353) and (hState = 331)) or
								((vState = 353) and (hState = 372)) or
								((vState = 353) and (hState = 382)) or
								((vState = 353) and (hState = 385)) or
								((vState = 353) and (hState = 439)) or
								((vState = 353) and (hState = 447)) or
								((vState = 353) and (hState = 448)) or
								((vState = 353) and (hState = 476)) or
								((vState = 353) and (hState = 477)) or
								((vState = 353) and (hState = 487)) or
								((vState = 353) and (hState = 488)) or
								((vState = 353) and (hState = 501)) or
								((vState = 353) and (hState = 507)) or
								((vState = 353) and (hState = 513)) or
								((vState = 353) and (hState = 514)) or
								((vState = 353) and (hState = 525)) or
								((vState = 353) and (hState = 526)) or
								((vState = 353) and (hState = 527)) or
								((vState = 353) and (hState = 541)) or
								((vState = 353) and (hState = 558)) or
								((vState = 353) and (hState = 559)) or
								((vState = 353) and (hState = 560)) or
								((vState = 353) and (hState = 561)) or
								((vState = 353) and (hState = 562)) or
								((vState = 353) and (hState = 563)) or
								((vState = 353) and (hState = 572)) or
								((vState = 353) and (hState = 573)) or
								((vState = 353) and (hState = 574)) or
								((vState = 353) and (hState = 575)) or
								((vState = 353) and (hState = 576)) or
								((vState = 353) and (hState = 577)) or
								((vState = 354) and (hState = 293)) or
								((vState = 354) and (hState = 294)) or
								((vState = 354) and (hState = 299)) or
								((vState = 354) and (hState = 300)) or
								((vState = 354) and (hState = 301)) or
								((vState = 354) and (hState = 308)) or
								((vState = 354) and (hState = 314)) or
								((vState = 354) and (hState = 328)) or
								((vState = 354) and (hState = 329)) or
								((vState = 354) and (hState = 330)) or
								((vState = 354) and (hState = 383)) or
								((vState = 354) and (hState = 384)) or
								((vState = 354) and (hState = 401)) or
								((vState = 354) and (hState = 402)) or
								((vState = 354) and (hState = 403)) or
								((vState = 354) and (hState = 418)) or
								((vState = 354) and (hState = 439)) or
								((vState = 354) and (hState = 448)) or
								((vState = 354) and (hState = 449)) or
								((vState = 354) and (hState = 450)) or
								((vState = 354) and (hState = 451)) or
								((vState = 354) and (hState = 452)) or
								((vState = 354) and (hState = 453)) or
								((vState = 354) and (hState = 454)) or
								((vState = 354) and (hState = 479)) or
								((vState = 354) and (hState = 480)) or
								((vState = 354) and (hState = 486)) or
								((vState = 354) and (hState = 487)) or
								((vState = 354) and (hState = 501)) or
								((vState = 354) and (hState = 502)) or
								((vState = 354) and (hState = 503)) or
								((vState = 354) and (hState = 507)) or
								((vState = 354) and (hState = 511)) or
								((vState = 354) and (hState = 512)) or
								((vState = 354) and (hState = 521)) or
								((vState = 354) and (hState = 522)) or
								((vState = 354) and (hState = 523)) or
								((vState = 354) and (hState = 524)) or
								((vState = 354) and (hState = 540)) or
								((vState = 354) and (hState = 541)) or
								((vState = 354) and (hState = 561)) or
								((vState = 354) and (hState = 562)) or
								((vState = 354) and (hState = 563)) or
								((vState = 354) and (hState = 564)) or
								((vState = 354) and (hState = 574)) or
								((vState = 354) and (hState = 575)) or
								((vState = 354) and (hState = 576)) or
								((vState = 354) and (hState = 577)) or
								((vState = 354) and (hState = 578)) or
								((vState = 354) and (hState = 579)) or
								((vState = 355) and (hState = 293)) or
								((vState = 355) and (hState = 294)) or
								((vState = 355) and (hState = 308)) or
								((vState = 355) and (hState = 315)) or
								((vState = 355) and (hState = 324)) or
								((vState = 355) and (hState = 325)) or
								((vState = 355) and (hState = 326)) or
								((vState = 355) and (hState = 327)) or
								((vState = 355) and (hState = 328)) or
								((vState = 355) and (hState = 329)) or
								((vState = 355) and (hState = 330)) or
								((vState = 355) and (hState = 383)) or
								((vState = 355) and (hState = 384)) or
								((vState = 355) and (hState = 401)) or
								((vState = 355) and (hState = 402)) or
								((vState = 355) and (hState = 413)) or
								((vState = 355) and (hState = 417)) or
								((vState = 355) and (hState = 448)) or
								((vState = 355) and (hState = 452)) or
								((vState = 355) and (hState = 453)) or
								((vState = 355) and (hState = 454)) or
								((vState = 355) and (hState = 455)) or
								((vState = 355) and (hState = 482)) or
								((vState = 355) and (hState = 486)) or
								((vState = 355) and (hState = 505)) or
								((vState = 355) and (hState = 506)) or
								((vState = 355) and (hState = 507)) or
								((vState = 355) and (hState = 508)) or
								((vState = 355) and (hState = 521)) or
								((vState = 355) and (hState = 522)) or
								((vState = 355) and (hState = 523)) or
								((vState = 355) and (hState = 524)) or
								((vState = 355) and (hState = 540)) or
								((vState = 355) and (hState = 541)) or
								((vState = 355) and (hState = 563)) or
								((vState = 355) and (hState = 564)) or
								((vState = 355) and (hState = 565)) or
								((vState = 355) and (hState = 578)) or
								((vState = 355) and (hState = 579)) or
								((vState = 355) and (hState = 580)) or
								((vState = 355) and (hState = 581)) or
								((vState = 355) and (hState = 582)) or
								((vState = 355) and (hState = 583)) or
								((vState = 356) and (hState = 293)) or
								((vState = 356) and (hState = 294)) or
								((vState = 356) and (hState = 308)) or
								((vState = 356) and (hState = 324)) or
								((vState = 356) and (hState = 325)) or
								((vState = 356) and (hState = 329)) or
								((vState = 356) and (hState = 330)) or
								((vState = 356) and (hState = 337)) or
								((vState = 356) and (hState = 383)) or
								((vState = 356) and (hState = 384)) or
								((vState = 356) and (hState = 401)) or
								((vState = 356) and (hState = 402)) or
								((vState = 356) and (hState = 448)) or
								((vState = 356) and (hState = 486)) or
								((vState = 356) and (hState = 505)) or
								((vState = 356) and (hState = 506)) or
								((vState = 356) and (hState = 507)) or
								((vState = 356) and (hState = 508)) or
								((vState = 356) and (hState = 563)) or
								((vState = 356) and (hState = 564)) or
								((vState = 356) and (hState = 565)) or
								((vState = 356) and (hState = 566)) or
								((vState = 356) and (hState = 581)) or
								((vState = 356) and (hState = 582)) or
								((vState = 356) and (hState = 583)) or
								((vState = 357) and (hState = 262)) or
								((vState = 357) and (hState = 293)) or
								((vState = 357) and (hState = 294)) or
								((vState = 357) and (hState = 308)) or
								((vState = 357) and (hState = 318)) or
								((vState = 357) and (hState = 321)) or
								((vState = 357) and (hState = 322)) or
								((vState = 357) and (hState = 323)) or
								((vState = 357) and (hState = 324)) or
								((vState = 357) and (hState = 329)) or
								((vState = 357) and (hState = 330)) or
								((vState = 357) and (hState = 336)) or
								((vState = 357) and (hState = 337)) or
								((vState = 357) and (hState = 383)) or
								((vState = 357) and (hState = 384)) or
								((vState = 357) and (hState = 401)) or
								((vState = 357) and (hState = 438)) or
								((vState = 357) and (hState = 448)) or
								((vState = 357) and (hState = 504)) or
								((vState = 357) and (hState = 505)) or
								((vState = 357) and (hState = 506)) or
								((vState = 357) and (hState = 507)) or
								((vState = 357) and (hState = 508)) or
								((vState = 357) and (hState = 545)) or
								((vState = 357) and (hState = 546)) or
								((vState = 357) and (hState = 563)) or
								((vState = 357) and (hState = 564)) or
								((vState = 357) and (hState = 565)) or
								((vState = 357) and (hState = 566)) or
								((vState = 357) and (hState = 567)) or
								((vState = 357) and (hState = 583)) or
								((vState = 357) and (hState = 584)) or
								((vState = 357) and (hState = 585)) or
								((vState = 357) and (hState = 590)) or
								((vState = 358) and (hState = 262)) or
								((vState = 358) and (hState = 292)) or
								((vState = 358) and (hState = 293)) or
								((vState = 358) and (hState = 294)) or
								((vState = 358) and (hState = 295)) or
								((vState = 358) and (hState = 296)) or
								((vState = 358) and (hState = 308)) or
								((vState = 358) and (hState = 318)) or
								((vState = 358) and (hState = 319)) or
								((vState = 358) and (hState = 320)) or
								((vState = 358) and (hState = 321)) or
								((vState = 358) and (hState = 322)) or
								((vState = 358) and (hState = 323)) or
								((vState = 358) and (hState = 329)) or
								((vState = 358) and (hState = 330)) or
								((vState = 358) and (hState = 336)) or
								((vState = 358) and (hState = 337)) or
								((vState = 358) and (hState = 383)) or
								((vState = 358) and (hState = 384)) or
								((vState = 358) and (hState = 401)) or
								((vState = 358) and (hState = 438)) or
								((vState = 358) and (hState = 448)) or
								((vState = 358) and (hState = 449)) or
								((vState = 358) and (hState = 450)) or
								((vState = 358) and (hState = 498)) or
								((vState = 358) and (hState = 503)) or
								((vState = 358) and (hState = 504)) or
								((vState = 358) and (hState = 511)) or
								((vState = 358) and (hState = 512)) or
								((vState = 358) and (hState = 513)) or
								((vState = 358) and (hState = 514)) or
								((vState = 358) and (hState = 515)) or
								((vState = 358) and (hState = 527)) or
								((vState = 358) and (hState = 537)) or
								((vState = 358) and (hState = 546)) or
								((vState = 358) and (hState = 556)) or
								((vState = 358) and (hState = 562)) or
								((vState = 358) and (hState = 563)) or
								((vState = 358) and (hState = 568)) or
								((vState = 358) and (hState = 585)) or
								((vState = 358) and (hState = 586)) or
								((vState = 358) and (hState = 587)) or
								((vState = 358) and (hState = 588)) or
								((vState = 358) and (hState = 589)) or
								((vState = 358) and (hState = 590)) or
								((vState = 359) and (hState = 292)) or
								((vState = 359) and (hState = 293)) or
								((vState = 359) and (hState = 294)) or
								((vState = 359) and (hState = 295)) or
								((vState = 359) and (hState = 304)) or
								((vState = 359) and (hState = 308)) or
								((vState = 359) and (hState = 318)) or
								((vState = 359) and (hState = 319)) or
								((vState = 359) and (hState = 320)) or
								((vState = 359) and (hState = 321)) or
								((vState = 359) and (hState = 322)) or
								((vState = 359) and (hState = 329)) or
								((vState = 359) and (hState = 330)) or
								((vState = 359) and (hState = 336)) or
								((vState = 359) and (hState = 344)) or
								((vState = 359) and (hState = 345)) or
								((vState = 359) and (hState = 346)) or
								((vState = 359) and (hState = 377)) or
								((vState = 359) and (hState = 383)) or
								((vState = 359) and (hState = 384)) or
								((vState = 359) and (hState = 400)) or
								((vState = 359) and (hState = 401)) or
								((vState = 359) and (hState = 434)) or
								((vState = 359) and (hState = 435)) or
								((vState = 359) and (hState = 436)) or
								((vState = 359) and (hState = 437)) or
								((vState = 359) and (hState = 438)) or
								((vState = 359) and (hState = 439)) or
								((vState = 359) and (hState = 440)) or
								((vState = 359) and (hState = 441)) or
								((vState = 359) and (hState = 442)) or
								((vState = 359) and (hState = 443)) or
								((vState = 359) and (hState = 444)) or
								((vState = 359) and (hState = 448)) or
								((vState = 359) and (hState = 449)) or
								((vState = 359) and (hState = 450)) or
								((vState = 359) and (hState = 465)) or
								((vState = 359) and (hState = 466)) or
								((vState = 359) and (hState = 490)) or
								((vState = 359) and (hState = 491)) or
								((vState = 359) and (hState = 492)) or
								((vState = 359) and (hState = 493)) or
								((vState = 359) and (hState = 494)) or
								((vState = 359) and (hState = 495)) or
								((vState = 359) and (hState = 496)) or
								((vState = 359) and (hState = 497)) or
								((vState = 359) and (hState = 498)) or
								((vState = 359) and (hState = 499)) or
								((vState = 359) and (hState = 500)) or
								((vState = 359) and (hState = 501)) or
								((vState = 359) and (hState = 502)) or
								((vState = 359) and (hState = 503)) or
								((vState = 359) and (hState = 512)) or
								((vState = 359) and (hState = 513)) or
								((vState = 359) and (hState = 514)) or
								((vState = 359) and (hState = 528)) or
								((vState = 359) and (hState = 537)) or
								((vState = 359) and (hState = 546)) or
								((vState = 359) and (hState = 556)) or
								((vState = 359) and (hState = 562)) or
								((vState = 359) and (hState = 568)) or
								((vState = 359) and (hState = 569)) or
								((vState = 359) and (hState = 585)) or
								((vState = 359) and (hState = 586)) or
								((vState = 359) and (hState = 587)) or
								((vState = 359) and (hState = 588)) or
								((vState = 359) and (hState = 589)) or
								((vState = 359) and (hState = 590)) or
								((vState = 359) and (hState = 591)) or
								((vState = 359) and (hState = 592)) or
								((vState = 359) and (hState = 593)) or
								((vState = 360) and (hState = 261)) or
								((vState = 360) and (hState = 292)) or
								((vState = 360) and (hState = 293)) or
								((vState = 360) and (hState = 294)) or
								((vState = 360) and (hState = 309)) or
								((vState = 360) and (hState = 317)) or
								((vState = 360) and (hState = 318)) or
								((vState = 360) and (hState = 319)) or
								((vState = 360) and (hState = 320)) or
								((vState = 360) and (hState = 321)) or
								((vState = 360) and (hState = 322)) or
								((vState = 360) and (hState = 331)) or
								((vState = 360) and (hState = 336)) or
								((vState = 360) and (hState = 350)) or
								((vState = 360) and (hState = 351)) or
								((vState = 360) and (hState = 352)) or
								((vState = 360) and (hState = 378)) or
								((vState = 360) and (hState = 383)) or
								((vState = 360) and (hState = 384)) or
								((vState = 360) and (hState = 400)) or
								((vState = 360) and (hState = 431)) or
								((vState = 360) and (hState = 432)) or
								((vState = 360) and (hState = 437)) or
								((vState = 360) and (hState = 447)) or
								((vState = 360) and (hState = 448)) or
								((vState = 360) and (hState = 449)) or
								((vState = 360) and (hState = 450)) or
								((vState = 360) and (hState = 451)) or
								((vState = 360) and (hState = 452)) or
								((vState = 360) and (hState = 453)) or
								((vState = 360) and (hState = 469)) or
								((vState = 360) and (hState = 470)) or
								((vState = 360) and (hState = 482)) or
								((vState = 360) and (hState = 496)) or
								((vState = 360) and (hState = 497)) or
								((vState = 360) and (hState = 514)) or
								((vState = 360) and (hState = 529)) or
								((vState = 360) and (hState = 536)) or
								((vState = 360) and (hState = 547)) or
								((vState = 360) and (hState = 556)) or
								((vState = 360) and (hState = 562)) or
								((vState = 360) and (hState = 588)) or
								((vState = 360) and (hState = 589)) or
								((vState = 360) and (hState = 590)) or
								((vState = 360) and (hState = 591)) or
								((vState = 360) and (hState = 592)) or
								((vState = 360) and (hState = 593)) or
								((vState = 360) and (hState = 594)) or
								((vState = 360) and (hState = 595)) or
								((vState = 361) and (hState = 261)) or
								((vState = 361) and (hState = 292)) or
								((vState = 361) and (hState = 293)) or
								((vState = 361) and (hState = 294)) or
								((vState = 361) and (hState = 309)) or
								((vState = 361) and (hState = 316)) or
								((vState = 361) and (hState = 317)) or
								((vState = 361) and (hState = 318)) or
								((vState = 361) and (hState = 319)) or
								((vState = 361) and (hState = 331)) or
								((vState = 361) and (hState = 336)) or
								((vState = 361) and (hState = 358)) or
								((vState = 361) and (hState = 383)) or
								((vState = 361) and (hState = 384)) or
								((vState = 361) and (hState = 437)) or
								((vState = 361) and (hState = 447)) or
								((vState = 361) and (hState = 448)) or
								((vState = 361) and (hState = 449)) or
								((vState = 361) and (hState = 496)) or
								((vState = 361) and (hState = 562)) or
								((vState = 361) and (hState = 590)) or
								((vState = 361) and (hState = 594)) or
								((vState = 361) and (hState = 595)) or
								((vState = 361) and (hState = 596)) or
								((vState = 362) and (hState = 292)) or
								((vState = 362) and (hState = 293)) or
								((vState = 362) and (hState = 309)) or
								((vState = 362) and (hState = 317)) or
								((vState = 362) and (hState = 318)) or
								((vState = 362) and (hState = 326)) or
								((vState = 362) and (hState = 358)) or
								((vState = 362) and (hState = 437)) or
								((vState = 362) and (hState = 447)) or
								((vState = 362) and (hState = 448)) or
								((vState = 362) and (hState = 449)) or
								((vState = 362) and (hState = 481)) or
								((vState = 362) and (hState = 558)) or
								((vState = 362) and (hState = 562)) or
								((vState = 362) and (hState = 590)) or
								((vState = 362) and (hState = 599)) or
								((vState = 363) and (hState = 267)) or
								((vState = 363) and (hState = 291)) or
								((vState = 363) and (hState = 292)) or
								((vState = 363) and (hState = 308)) or
								((vState = 363) and (hState = 309)) or
								((vState = 363) and (hState = 326)) or
								((vState = 363) and (hState = 385)) or
								((vState = 363) and (hState = 397)) or
								((vState = 363) and (hState = 398)) or
								((vState = 363) and (hState = 449)) or
								((vState = 363) and (hState = 480)) or
								((vState = 363) and (hState = 532)) or
								((vState = 363) and (hState = 559)) or
								((vState = 363) and (hState = 560)) or
								((vState = 363) and (hState = 561)) or
								((vState = 363) and (hState = 562)) or
								((vState = 363) and (hState = 590)) or
								((vState = 364) and (hState = 260)) or
								((vState = 364) and (hState = 267)) or
								((vState = 364) and (hState = 291)) or
								((vState = 364) and (hState = 292)) or
								((vState = 364) and (hState = 308)) or
								((vState = 364) and (hState = 309)) or
								((vState = 364) and (hState = 310)) or
								((vState = 364) and (hState = 311)) or
								((vState = 364) and (hState = 326)) or
								((vState = 364) and (hState = 327)) or
								((vState = 364) and (hState = 333)) or
								((vState = 364) and (hState = 334)) or
								((vState = 364) and (hState = 335)) or
								((vState = 364) and (hState = 367)) or
								((vState = 364) and (hState = 368)) or
								((vState = 364) and (hState = 369)) or
								((vState = 364) and (hState = 370)) or
								((vState = 364) and (hState = 371)) or
								((vState = 364) and (hState = 381)) or
								((vState = 364) and (hState = 382)) or
								((vState = 364) and (hState = 385)) or
								((vState = 364) and (hState = 396)) or
								((vState = 364) and (hState = 397)) or
								((vState = 364) and (hState = 418)) or
								((vState = 364) and (hState = 419)) or
								((vState = 364) and (hState = 445)) or
								((vState = 364) and (hState = 449)) or
								((vState = 364) and (hState = 464)) or
								((vState = 364) and (hState = 480)) or
								((vState = 364) and (hState = 532)) or
								((vState = 364) and (hState = 533)) or
								((vState = 364) and (hState = 534)) or
								((vState = 364) and (hState = 553)) or
								((vState = 364) and (hState = 560)) or
								((vState = 364) and (hState = 561)) or
								((vState = 364) and (hState = 562)) or
								((vState = 364) and (hState = 590)) or
								((vState = 365) and (hState = 260)) or
								((vState = 365) and (hState = 261)) or
								((vState = 365) and (hState = 262)) or
								((vState = 365) and (hState = 267)) or
								((vState = 365) and (hState = 308)) or
								((vState = 365) and (hState = 309)) or
								((vState = 365) and (hState = 310)) or
								((vState = 365) and (hState = 311)) or
								((vState = 365) and (hState = 315)) or
								((vState = 365) and (hState = 325)) or
								((vState = 365) and (hState = 330)) or
								((vState = 365) and (hState = 331)) or
								((vState = 365) and (hState = 332)) or
								((vState = 365) and (hState = 333)) or
								((vState = 365) and (hState = 334)) or
								((vState = 365) and (hState = 335)) or
								((vState = 365) and (hState = 368)) or
								((vState = 365) and (hState = 369)) or
								((vState = 365) and (hState = 370)) or
								((vState = 365) and (hState = 371)) or
								((vState = 365) and (hState = 382)) or
								((vState = 365) and (hState = 385)) or
								((vState = 365) and (hState = 396)) or
								((vState = 365) and (hState = 397)) or
								((vState = 365) and (hState = 415)) or
								((vState = 365) and (hState = 416)) or
								((vState = 365) and (hState = 444)) or
								((vState = 365) and (hState = 449)) or
								((vState = 365) and (hState = 466)) or
								((vState = 365) and (hState = 480)) or
								((vState = 365) and (hState = 523)) or
								((vState = 365) and (hState = 532)) or
								((vState = 365) and (hState = 533)) or
								((vState = 365) and (hState = 534)) or
								((vState = 365) and (hState = 561)) or
								((vState = 365) and (hState = 562)) or
								((vState = 365) and (hState = 563)) or
								((vState = 365) and (hState = 564)) or
								((vState = 365) and (hState = 577)) or
								((vState = 365) and (hState = 590)) or
								((vState = 366) and (hState = 260)) or
								((vState = 366) and (hState = 267)) or
								((vState = 366) and (hState = 308)) or
								((vState = 366) and (hState = 309)) or
								((vState = 366) and (hState = 310)) or
								((vState = 366) and (hState = 311)) or
								((vState = 366) and (hState = 312)) or
								((vState = 366) and (hState = 313)) or
								((vState = 366) and (hState = 325)) or
								((vState = 366) and (hState = 331)) or
								((vState = 366) and (hState = 332)) or
								((vState = 366) and (hState = 333)) or
								((vState = 366) and (hState = 334)) or
								((vState = 366) and (hState = 335)) or
								((vState = 366) and (hState = 368)) or
								((vState = 366) and (hState = 382)) or
								((vState = 366) and (hState = 383)) or
								((vState = 366) and (hState = 384)) or
								((vState = 366) and (hState = 385)) or
								((vState = 366) and (hState = 395)) or
								((vState = 366) and (hState = 396)) or
								((vState = 366) and (hState = 411)) or
								((vState = 366) and (hState = 412)) or
								((vState = 366) and (hState = 443)) or
								((vState = 366) and (hState = 449)) or
								((vState = 366) and (hState = 525)) or
								((vState = 366) and (hState = 532)) or
								((vState = 366) and (hState = 533)) or
								((vState = 366) and (hState = 534)) or
								((vState = 366) and (hState = 535)) or
								((vState = 366) and (hState = 557)) or
								((vState = 366) and (hState = 561)) or
								((vState = 366) and (hState = 562)) or
								((vState = 366) and (hState = 563)) or
								((vState = 366) and (hState = 564)) or
								((vState = 366) and (hState = 565)) or
								((vState = 367) and (hState = 267)) or
								((vState = 367) and (hState = 310)) or
								((vState = 367) and (hState = 311)) or
								((vState = 367) and (hState = 312)) or
								((vState = 367) and (hState = 313)) or
								((vState = 367) and (hState = 325)) or
								((vState = 367) and (hState = 334)) or
								((vState = 367) and (hState = 335)) or
								((vState = 367) and (hState = 384)) or
								((vState = 367) and (hState = 385)) or
								((vState = 367) and (hState = 395)) or
								((vState = 367) and (hState = 396)) or
								((vState = 367) and (hState = 449)) or
								((vState = 367) and (hState = 532)) or
								((vState = 367) and (hState = 561)) or
								((vState = 367) and (hState = 565)) or
								((vState = 367) and (hState = 566)) or
								((vState = 368) and (hState = 257)) or
								((vState = 368) and (hState = 258)) or
								((vState = 368) and (hState = 267)) or
								((vState = 368) and (hState = 310)) or
								((vState = 368) and (hState = 311)) or
								((vState = 368) and (hState = 312)) or
								((vState = 368) and (hState = 313)) or
								((vState = 368) and (hState = 334)) or
								((vState = 368) and (hState = 335)) or
								((vState = 368) and (hState = 385)) or
								((vState = 368) and (hState = 386)) or
								((vState = 368) and (hState = 387)) or
								((vState = 368) and (hState = 394)) or
								((vState = 368) and (hState = 395)) or
								((vState = 368) and (hState = 449)) or
								((vState = 368) and (hState = 560)) or
								((vState = 368) and (hState = 566)) or
								((vState = 368) and (hState = 567)) or
								((vState = 368) and (hState = 568)) or
								((vState = 369) and (hState = 256)) or
								((vState = 369) and (hState = 257)) or
								((vState = 369) and (hState = 258)) or
								((vState = 369) and (hState = 267)) or
								((vState = 369) and (hState = 304)) or
								((vState = 369) and (hState = 310)) or
								((vState = 369) and (hState = 311)) or
								((vState = 369) and (hState = 312)) or
								((vState = 369) and (hState = 313)) or
								((vState = 369) and (hState = 334)) or
								((vState = 369) and (hState = 335)) or
								((vState = 369) and (hState = 357)) or
								((vState = 369) and (hState = 363)) or
								((vState = 369) and (hState = 385)) or
								((vState = 369) and (hState = 386)) or
								((vState = 369) and (hState = 387)) or
								((vState = 369) and (hState = 392)) or
								((vState = 369) and (hState = 393)) or
								((vState = 369) and (hState = 394)) or
								((vState = 369) and (hState = 395)) or
								((vState = 369) and (hState = 402)) or
								((vState = 369) and (hState = 403)) or
								((vState = 369) and (hState = 434)) or
								((vState = 369) and (hState = 449)) or
								((vState = 369) and (hState = 470)) or
								((vState = 369) and (hState = 492)) or
								((vState = 369) and (hState = 529)) or
								((vState = 369) and (hState = 530)) or
								((vState = 369) and (hState = 531)) or
								((vState = 369) and (hState = 560)) or
								((vState = 369) and (hState = 561)) or
								((vState = 369) and (hState = 566)) or
								((vState = 369) and (hState = 567)) or
								((vState = 369) and (hState = 568)) or
								((vState = 369) and (hState = 569)) or
								((vState = 369) and (hState = 570)) or
								((vState = 369) and (hState = 589)) or
								((vState = 370) and (hState = 267)) or
								((vState = 370) and (hState = 309)) or
								((vState = 370) and (hState = 310)) or
								((vState = 370) and (hState = 311)) or
								((vState = 370) and (hState = 312)) or
								((vState = 370) and (hState = 313)) or
								((vState = 370) and (hState = 326)) or
								((vState = 370) and (hState = 334)) or
								((vState = 370) and (hState = 335)) or
								((vState = 370) and (hState = 336)) or
								((vState = 370) and (hState = 337)) or
								((vState = 370) and (hState = 357)) or
								((vState = 370) and (hState = 361)) or
								((vState = 370) and (hState = 386)) or
								((vState = 370) and (hState = 387)) or
								((vState = 370) and (hState = 392)) or
								((vState = 370) and (hState = 393)) or
								((vState = 370) and (hState = 394)) or
								((vState = 370) and (hState = 395)) or
								((vState = 370) and (hState = 399)) or
								((vState = 370) and (hState = 400)) or
								((vState = 370) and (hState = 434)) or
								((vState = 370) and (hState = 449)) or
								((vState = 370) and (hState = 471)) or
								((vState = 370) and (hState = 476)) or
								((vState = 370) and (hState = 540)) or
								((vState = 370) and (hState = 561)) or
								((vState = 370) and (hState = 562)) or
								((vState = 370) and (hState = 567)) or
								((vState = 370) and (hState = 568)) or
								((vState = 370) and (hState = 572)) or
								((vState = 370) and (hState = 583)) or
								((vState = 370) and (hState = 589)) or
								((vState = 371) and (hState = 251)) or
								((vState = 371) and (hState = 252)) or
								((vState = 371) and (hState = 267)) or
								((vState = 371) and (hState = 313)) or
								((vState = 371) and (hState = 314)) or
								((vState = 371) and (hState = 326)) or
								((vState = 371) and (hState = 327)) or
								((vState = 371) and (hState = 331)) or
								((vState = 371) and (hState = 332)) or
								((vState = 371) and (hState = 333)) or
								((vState = 371) and (hState = 334)) or
								((vState = 371) and (hState = 335)) or
								((vState = 371) and (hState = 336)) or
								((vState = 371) and (hState = 337)) or
								((vState = 371) and (hState = 338)) or
								((vState = 371) and (hState = 357)) or
								((vState = 371) and (hState = 358)) or
								((vState = 371) and (hState = 386)) or
								((vState = 371) and (hState = 387)) or
								((vState = 371) and (hState = 388)) or
								((vState = 371) and (hState = 391)) or
								((vState = 371) and (hState = 392)) or
								((vState = 371) and (hState = 393)) or
								((vState = 371) and (hState = 394)) or
								((vState = 371) and (hState = 395)) or
								((vState = 371) and (hState = 396)) or
								((vState = 371) and (hState = 431)) or
								((vState = 371) and (hState = 432)) or
								((vState = 371) and (hState = 433)) or
								((vState = 371) and (hState = 434)) or
								((vState = 371) and (hState = 439)) or
								((vState = 371) and (hState = 449)) or
								((vState = 371) and (hState = 474)) or
								((vState = 371) and (hState = 475)) or
								((vState = 371) and (hState = 491)) or
								((vState = 371) and (hState = 514)) or
								((vState = 371) and (hState = 541)) or
								((vState = 371) and (hState = 561)) or
								((vState = 371) and (hState = 562)) or
								((vState = 371) and (hState = 563)) or
								((vState = 371) and (hState = 567)) or
								((vState = 371) and (hState = 568)) or
								((vState = 371) and (hState = 574)) or
								((vState = 371) and (hState = 584)) or
								((vState = 371) and (hState = 589)) or
								((vState = 372) and (hState = 267)) or
								((vState = 372) and (hState = 313)) or
								((vState = 372) and (hState = 314)) or
								((vState = 372) and (hState = 326)) or
								((vState = 372) and (hState = 327)) or
								((vState = 372) and (hState = 328)) or
								((vState = 372) and (hState = 336)) or
								((vState = 372) and (hState = 357)) or
								((vState = 372) and (hState = 388)) or
								((vState = 372) and (hState = 391)) or
								((vState = 372) and (hState = 392)) or
								((vState = 372) and (hState = 393)) or
								((vState = 372) and (hState = 433)) or
								((vState = 372) and (hState = 434)) or
								((vState = 372) and (hState = 439)) or
								((vState = 372) and (hState = 449)) or
								((vState = 372) and (hState = 475)) or
								((vState = 372) and (hState = 561)) or
								((vState = 372) and (hState = 567)) or
								((vState = 372) and (hState = 568)) or
								((vState = 372) and (hState = 589)) or
								((vState = 373) and (hState = 257)) or
								((vState = 373) and (hState = 267)) or
								((vState = 373) and (hState = 288)) or
								((vState = 373) and (hState = 313)) or
								((vState = 373) and (hState = 314)) or
								((vState = 373) and (hState = 329)) or
								((vState = 373) and (hState = 336)) or
								((vState = 373) and (hState = 356)) or
								((vState = 373) and (hState = 379)) or
								((vState = 373) and (hState = 388)) or
								((vState = 373) and (hState = 389)) or
								((vState = 373) and (hState = 390)) or
								((vState = 373) and (hState = 391)) or
								((vState = 373) and (hState = 392)) or
								((vState = 373) and (hState = 433)) or
								((vState = 373) and (hState = 434)) or
								((vState = 373) and (hState = 435)) or
								((vState = 373) and (hState = 436)) or
								((vState = 373) and (hState = 437)) or
								((vState = 373) and (hState = 438)) or
								((vState = 373) and (hState = 439)) or
								((vState = 373) and (hState = 449)) or
								((vState = 373) and (hState = 475)) or
								((vState = 373) and (hState = 490)) or
								((vState = 373) and (hState = 567)) or
								((vState = 373) and (hState = 568)) or
								((vState = 373) and (hState = 569)) or
								((vState = 373) and (hState = 589)) or
								((vState = 374) and (hState = 257)) or
								((vState = 374) and (hState = 267)) or
								((vState = 374) and (hState = 288)) or
								((vState = 374) and (hState = 297)) or
								((vState = 374) and (hState = 304)) or
								((vState = 374) and (hState = 313)) or
								((vState = 374) and (hState = 314)) or
								((vState = 374) and (hState = 315)) or
								((vState = 374) and (hState = 319)) or
								((vState = 374) and (hState = 320)) or
								((vState = 374) and (hState = 321)) or
								((vState = 374) and (hState = 322)) or
								((vState = 374) and (hState = 329)) or
								((vState = 374) and (hState = 336)) or
								((vState = 374) and (hState = 354)) or
								((vState = 374) and (hState = 355)) or
								((vState = 374) and (hState = 356)) or
								((vState = 374) and (hState = 379)) or
								((vState = 374) and (hState = 388)) or
								((vState = 374) and (hState = 389)) or
								((vState = 374) and (hState = 390)) or
								((vState = 374) and (hState = 391)) or
								((vState = 374) and (hState = 392)) or
								((vState = 374) and (hState = 433)) or
								((vState = 374) and (hState = 434)) or
								((vState = 374) and (hState = 435)) or
								((vState = 374) and (hState = 436)) or
								((vState = 374) and (hState = 437)) or
								((vState = 374) and (hState = 438)) or
								((vState = 374) and (hState = 439)) or
								((vState = 374) and (hState = 440)) or
								((vState = 374) and (hState = 449)) or
								((vState = 374) and (hState = 475)) or
								((vState = 374) and (hState = 476)) or
								((vState = 374) and (hState = 490)) or
								((vState = 374) and (hState = 496)) or
								((vState = 374) and (hState = 497)) or
								((vState = 374) and (hState = 498)) or
								((vState = 374) and (hState = 518)) or
								((vState = 374) and (hState = 519)) or
								((vState = 374) and (hState = 561)) or
								((vState = 374) and (hState = 567)) or
								((vState = 374) and (hState = 568)) or
								((vState = 374) and (hState = 569)) or
								((vState = 374) and (hState = 570)) or
								((vState = 374) and (hState = 578)) or
								((vState = 374) and (hState = 579)) or
								((vState = 374) and (hState = 588)) or
								((vState = 374) and (hState = 589)) or
								((vState = 375) and (hState = 246)) or
								((vState = 375) and (hState = 257)) or
								((vState = 375) and (hState = 267)) or
								((vState = 375) and (hState = 288)) or
								((vState = 375) and (hState = 304)) or
								((vState = 375) and (hState = 313)) or
								((vState = 375) and (hState = 314)) or
								((vState = 375) and (hState = 315)) or
								((vState = 375) and (hState = 316)) or
								((vState = 375) and (hState = 330)) or
								((vState = 375) and (hState = 331)) or
								((vState = 375) and (hState = 332)) or
								((vState = 375) and (hState = 344)) or
								((vState = 375) and (hState = 345)) or
								((vState = 375) and (hState = 351)) or
								((vState = 375) and (hState = 352)) or
								((vState = 375) and (hState = 356)) or
								((vState = 375) and (hState = 379)) or
								((vState = 375) and (hState = 388)) or
								((vState = 375) and (hState = 389)) or
								((vState = 375) and (hState = 390)) or
								((vState = 375) and (hState = 391)) or
								((vState = 375) and (hState = 433)) or
								((vState = 375) and (hState = 434)) or
								((vState = 375) and (hState = 435)) or
								((vState = 375) and (hState = 442)) or
								((vState = 375) and (hState = 443)) or
								((vState = 375) and (hState = 444)) or
								((vState = 375) and (hState = 449)) or
								((vState = 375) and (hState = 474)) or
								((vState = 375) and (hState = 489)) or
								((vState = 375) and (hState = 490)) or
								((vState = 375) and (hState = 491)) or
								((vState = 375) and (hState = 492)) or
								((vState = 375) and (hState = 493)) or
								((vState = 375) and (hState = 545)) or
								((vState = 375) and (hState = 562)) or
								((vState = 375) and (hState = 568)) or
								((vState = 375) and (hState = 569)) or
								((vState = 375) and (hState = 570)) or
								((vState = 375) and (hState = 571)) or
								((vState = 375) and (hState = 572)) or
								((vState = 375) and (hState = 589)) or
								((vState = 375) and (hState = 599)) or
								((vState = 376) and (hState = 244)) or
								((vState = 376) and (hState = 257)) or
								((vState = 376) and (hState = 261)) or
								((vState = 376) and (hState = 262)) or
								((vState = 376) and (hState = 263)) or
								((vState = 376) and (hState = 293)) or
								((vState = 376) and (hState = 304)) or
								((vState = 376) and (hState = 305)) or
								((vState = 376) and (hState = 306)) or
								((vState = 376) and (hState = 307)) or
								((vState = 376) and (hState = 308)) or
								((vState = 376) and (hState = 309)) or
								((vState = 376) and (hState = 310)) or
								((vState = 376) and (hState = 315)) or
								((vState = 376) and (hState = 316)) or
								((vState = 376) and (hState = 331)) or
								((vState = 376) and (hState = 332)) or
								((vState = 376) and (hState = 346)) or
								((vState = 376) and (hState = 347)) or
								((vState = 376) and (hState = 348)) or
								((vState = 376) and (hState = 349)) or
								((vState = 376) and (hState = 350)) or
								((vState = 376) and (hState = 356)) or
								((vState = 376) and (hState = 388)) or
								((vState = 376) and (hState = 389)) or
								((vState = 376) and (hState = 390)) or
								((vState = 376) and (hState = 391)) or
								((vState = 376) and (hState = 432)) or
								((vState = 376) and (hState = 433)) or
								((vState = 376) and (hState = 434)) or
								((vState = 376) and (hState = 446)) or
								((vState = 376) and (hState = 447)) or
								((vState = 376) and (hState = 448)) or
								((vState = 376) and (hState = 449)) or
								((vState = 376) and (hState = 450)) or
								((vState = 376) and (hState = 474)) or
								((vState = 376) and (hState = 489)) or
								((vState = 376) and (hState = 490)) or
								((vState = 376) and (hState = 491)) or
								((vState = 376) and (hState = 501)) or
								((vState = 376) and (hState = 523)) or
								((vState = 376) and (hState = 545)) or
								((vState = 376) and (hState = 563)) or
								((vState = 376) and (hState = 571)) or
								((vState = 376) and (hState = 572)) or
								((vState = 376) and (hState = 573)) or
								((vState = 376) and (hState = 584)) or
								((vState = 376) and (hState = 589)) or
								((vState = 376) and (hState = 590)) or
								((vState = 377) and (hState = 257)) or
								((vState = 377) and (hState = 258)) or
								((vState = 377) and (hState = 293)) or
								((vState = 377) and (hState = 304)) or
								((vState = 377) and (hState = 331)) or
								((vState = 377) and (hState = 332)) or
								((vState = 377) and (hState = 346)) or
								((vState = 377) and (hState = 347)) or
								((vState = 377) and (hState = 348)) or
								((vState = 377) and (hState = 349)) or
								((vState = 377) and (hState = 350)) or
								((vState = 377) and (hState = 356)) or
								((vState = 377) and (hState = 387)) or
								((vState = 377) and (hState = 388)) or
								((vState = 377) and (hState = 389)) or
								((vState = 377) and (hState = 390)) or
								((vState = 377) and (hState = 391)) or
								((vState = 377) and (hState = 432)) or
								((vState = 377) and (hState = 433)) or
								((vState = 377) and (hState = 449)) or
								((vState = 377) and (hState = 450)) or
								((vState = 377) and (hState = 572)) or
								((vState = 377) and (hState = 573)) or
								((vState = 377) and (hState = 589)) or
								((vState = 377) and (hState = 590)) or
								((vState = 378) and (hState = 256)) or
								((vState = 378) and (hState = 287)) or
								((vState = 378) and (hState = 292)) or
								((vState = 378) and (hState = 293)) or
								((vState = 378) and (hState = 303)) or
								((vState = 378) and (hState = 331)) or
								((vState = 378) and (hState = 332)) or
								((vState = 378) and (hState = 350)) or
								((vState = 378) and (hState = 378)) or
								((vState = 378) and (hState = 386)) or
								((vState = 378) and (hState = 387)) or
								((vState = 378) and (hState = 388)) or
								((vState = 378) and (hState = 389)) or
								((vState = 378) and (hState = 390)) or
								((vState = 378) and (hState = 391)) or
								((vState = 378) and (hState = 392)) or
								((vState = 378) and (hState = 432)) or
								((vState = 378) and (hState = 481)) or
								((vState = 378) and (hState = 574)) or
								((vState = 378) and (hState = 575)) or
								((vState = 378) and (hState = 589)) or
								((vState = 378) and (hState = 590)) or
								((vState = 378) and (hState = 591)) or
								((vState = 379) and (hState = 255)) or
								((vState = 379) and (hState = 267)) or
								((vState = 379) and (hState = 287)) or
								((vState = 379) and (hState = 288)) or
								((vState = 379) and (hState = 289)) or
								((vState = 379) and (hState = 290)) or
								((vState = 379) and (hState = 291)) or
								((vState = 379) and (hState = 292)) or
								((vState = 379) and (hState = 303)) or
								((vState = 379) and (hState = 331)) or
								((vState = 379) and (hState = 332)) or
								((vState = 379) and (hState = 350)) or
								((vState = 379) and (hState = 378)) or
								((vState = 379) and (hState = 387)) or
								((vState = 379) and (hState = 388)) or
								((vState = 379) and (hState = 389)) or
								((vState = 379) and (hState = 390)) or
								((vState = 379) and (hState = 391)) or
								((vState = 379) and (hState = 393)) or
								((vState = 379) and (hState = 432)) or
								((vState = 379) and (hState = 452)) or
								((vState = 379) and (hState = 453)) or
								((vState = 379) and (hState = 481)) or
								((vState = 379) and (hState = 482)) or
								((vState = 379) and (hState = 483)) or
								((vState = 379) and (hState = 484)) or
								((vState = 379) and (hState = 485)) or
								((vState = 379) and (hState = 486)) or
								((vState = 379) and (hState = 527)) or
								((vState = 379) and (hState = 575)) or
								((vState = 379) and (hState = 576)) or
								((vState = 379) and (hState = 577)) or
								((vState = 379) and (hState = 591)) or
								((vState = 379) and (hState = 592)) or
								((vState = 379) and (hState = 593)) or
								((vState = 379) and (hState = 594)) or
								((vState = 379) and (hState = 595)) or
								((vState = 380) and (hState = 238)) or
								((vState = 380) and (hState = 250)) or
								((vState = 380) and (hState = 251)) or
								((vState = 380) and (hState = 255)) or
								((vState = 380) and (hState = 267)) or
								((vState = 380) and (hState = 268)) or
								((vState = 380) and (hState = 287)) or
								((vState = 380) and (hState = 288)) or
								((vState = 380) and (hState = 289)) or
								((vState = 380) and (hState = 290)) or
								((vState = 380) and (hState = 291)) or
								((vState = 380) and (hState = 292)) or
								((vState = 380) and (hState = 303)) or
								((vState = 380) and (hState = 318)) or
								((vState = 380) and (hState = 331)) or
								((vState = 380) and (hState = 332)) or
								((vState = 380) and (hState = 342)) or
								((vState = 380) and (hState = 351)) or
								((vState = 380) and (hState = 352)) or
								((vState = 380) and (hState = 353)) or
								((vState = 380) and (hState = 354)) or
								((vState = 380) and (hState = 355)) or
								((vState = 380) and (hState = 378)) or
								((vState = 380) and (hState = 384)) or
								((vState = 380) and (hState = 388)) or
								((vState = 380) and (hState = 389)) or
								((vState = 380) and (hState = 390)) or
								((vState = 380) and (hState = 394)) or
								((vState = 380) and (hState = 432)) or
								((vState = 380) and (hState = 453)) or
								((vState = 380) and (hState = 457)) or
								((vState = 380) and (hState = 458)) or
								((vState = 380) and (hState = 459)) or
								((vState = 380) and (hState = 476)) or
								((vState = 380) and (hState = 481)) or
								((vState = 380) and (hState = 482)) or
								((vState = 380) and (hState = 483)) or
								((vState = 380) and (hState = 484)) or
								((vState = 380) and (hState = 485)) or
								((vState = 380) and (hState = 486)) or
								((vState = 380) and (hState = 528)) or
								((vState = 380) and (hState = 529)) or
								((vState = 380) and (hState = 567)) or
								((vState = 380) and (hState = 576)) or
								((vState = 380) and (hState = 577)) or
								((vState = 380) and (hState = 578)) or
								((vState = 380) and (hState = 592)) or
								((vState = 380) and (hState = 593)) or
								((vState = 380) and (hState = 594)) or
								((vState = 380) and (hState = 595)) or
								((vState = 381) and (hState = 236)) or
								((vState = 381) and (hState = 237)) or
								((vState = 381) and (hState = 246)) or
								((vState = 381) and (hState = 247)) or
								((vState = 381) and (hState = 248)) or
								((vState = 381) and (hState = 255)) or
								((vState = 381) and (hState = 303)) or
								((vState = 381) and (hState = 331)) or
								((vState = 381) and (hState = 332)) or
								((vState = 381) and (hState = 333)) or
								((vState = 381) and (hState = 334)) or
								((vState = 381) and (hState = 339)) or
								((vState = 381) and (hState = 340)) or
								((vState = 381) and (hState = 341)) or
								((vState = 381) and (hState = 342)) or
								((vState = 381) and (hState = 351)) or
								((vState = 381) and (hState = 352)) or
								((vState = 381) and (hState = 353)) or
								((vState = 381) and (hState = 354)) or
								((vState = 381) and (hState = 355)) or
								((vState = 381) and (hState = 356)) or
								((vState = 381) and (hState = 357)) or
								((vState = 381) and (hState = 358)) or
								((vState = 381) and (hState = 359)) or
								((vState = 381) and (hState = 360)) or
								((vState = 381) and (hState = 361)) or
								((vState = 381) and (hState = 362)) or
								((vState = 381) and (hState = 363)) or
								((vState = 381) and (hState = 364)) or
								((vState = 381) and (hState = 365)) or
								((vState = 381) and (hState = 366)) or
								((vState = 381) and (hState = 367)) or
								((vState = 381) and (hState = 368)) or
								((vState = 381) and (hState = 369)) or
								((vState = 381) and (hState = 370)) or
								((vState = 381) and (hState = 371)) or
								((vState = 381) and (hState = 372)) or
								((vState = 381) and (hState = 373)) or
								((vState = 381) and (hState = 374)) or
								((vState = 381) and (hState = 388)) or
								((vState = 381) and (hState = 395)) or
								((vState = 381) and (hState = 460)) or
								((vState = 381) and (hState = 461)) or
								((vState = 381) and (hState = 462)) or
								((vState = 381) and (hState = 476)) or
								((vState = 381) and (hState = 477)) or
								((vState = 381) and (hState = 478)) or
								((vState = 381) and (hState = 485)) or
								((vState = 381) and (hState = 486)) or
								((vState = 381) and (hState = 506)) or
								((vState = 381) and (hState = 530)) or
								((vState = 381) and (hState = 568)) or
								((vState = 381) and (hState = 578)) or
								((vState = 381) and (hState = 579)) or
								((vState = 381) and (hState = 588)) or
								((vState = 381) and (hState = 593)) or
								((vState = 381) and (hState = 594)) or
								((vState = 381) and (hState = 595)) or
								((vState = 381) and (hState = 596)) or
								((vState = 382) and (hState = 255)) or
								((vState = 382) and (hState = 303)) or
								((vState = 382) and (hState = 331)) or
								((vState = 382) and (hState = 332)) or
								((vState = 382) and (hState = 333)) or
								((vState = 382) and (hState = 334)) or
								((vState = 382) and (hState = 338)) or
								((vState = 382) and (hState = 339)) or
								((vState = 382) and (hState = 340)) or
								((vState = 382) and (hState = 341)) or
								((vState = 382) and (hState = 342)) or
								((vState = 382) and (hState = 343)) or
								((vState = 382) and (hState = 355)) or
								((vState = 382) and (hState = 356)) or
								((vState = 382) and (hState = 357)) or
								((vState = 382) and (hState = 358)) or
								((vState = 382) and (hState = 383)) or
								((vState = 382) and (hState = 387)) or
								((vState = 382) and (hState = 388)) or
								((vState = 382) and (hState = 391)) or
								((vState = 382) and (hState = 396)) or
								((vState = 382) and (hState = 430)) or
								((vState = 382) and (hState = 476)) or
								((vState = 382) and (hState = 477)) or
								((vState = 382) and (hState = 478)) or
								((vState = 382) and (hState = 485)) or
								((vState = 382) and (hState = 486)) or
								((vState = 382) and (hState = 569)) or
								((vState = 382) and (hState = 579)) or
								((vState = 382) and (hState = 580)) or
								((vState = 382) and (hState = 588)) or
								((vState = 382) and (hState = 593)) or
								((vState = 382) and (hState = 597)) or
								((vState = 383) and (hState = 269)) or
								((vState = 383) and (hState = 319)) or
								((vState = 383) and (hState = 320)) or
								((vState = 383) and (hState = 330)) or
								((vState = 383) and (hState = 331)) or
								((vState = 383) and (hState = 332)) or
								((vState = 383) and (hState = 333)) or
								((vState = 383) and (hState = 334)) or
								((vState = 383) and (hState = 335)) or
								((vState = 383) and (hState = 336)) or
								((vState = 383) and (hState = 340)) or
								((vState = 383) and (hState = 341)) or
								((vState = 383) and (hState = 355)) or
								((vState = 383) and (hState = 356)) or
								((vState = 383) and (hState = 357)) or
								((vState = 383) and (hState = 358)) or
								((vState = 383) and (hState = 386)) or
								((vState = 383) and (hState = 387)) or
								((vState = 383) and (hState = 391)) or
								((vState = 383) and (hState = 405)) or
								((vState = 383) and (hState = 406)) or
								((vState = 383) and (hState = 429)) or
								((vState = 383) and (hState = 532)) or
								((vState = 383) and (hState = 533)) or
								((vState = 383) and (hState = 588)) or
								((vState = 384) and (hState = 232)) or
								((vState = 384) and (hState = 269)) or
								((vState = 384) and (hState = 270)) or
								((vState = 384) and (hState = 320)) or
								((vState = 384) and (hState = 330)) or
								((vState = 384) and (hState = 331)) or
								((vState = 384) and (hState = 332)) or
								((vState = 384) and (hState = 333)) or
								((vState = 384) and (hState = 334)) or
								((vState = 384) and (hState = 335)) or
								((vState = 384) and (hState = 336)) or
								((vState = 384) and (hState = 341)) or
								((vState = 384) and (hState = 357)) or
								((vState = 384) and (hState = 358)) or
								((vState = 384) and (hState = 385)) or
								((vState = 384) and (hState = 386)) or
								((vState = 384) and (hState = 387)) or
								((vState = 384) and (hState = 405)) or
								((vState = 384) and (hState = 406)) or
								((vState = 384) and (hState = 428)) or
								((vState = 384) and (hState = 429)) or
								((vState = 384) and (hState = 468)) or
								((vState = 384) and (hState = 469)) or
								((vState = 384) and (hState = 470)) or
								((vState = 384) and (hState = 471)) or
								((vState = 384) and (hState = 472)) or
								((vState = 384) and (hState = 473)) or
								((vState = 384) and (hState = 474)) or
								((vState = 384) and (hState = 532)) or
								((vState = 384) and (hState = 588)) or
								((vState = 385) and (hState = 231)) or
								((vState = 385) and (hState = 232)) or
								((vState = 385) and (hState = 236)) or
								((vState = 385) and (hState = 237)) or
								((vState = 385) and (hState = 238)) or
								((vState = 385) and (hState = 269)) or
								((vState = 385) and (hState = 270)) or
								((vState = 385) and (hState = 271)) or
								((vState = 385) and (hState = 281)) or
								((vState = 385) and (hState = 320)) or
								((vState = 385) and (hState = 330)) or
								((vState = 385) and (hState = 331)) or
								((vState = 385) and (hState = 332)) or
								((vState = 385) and (hState = 333)) or
								((vState = 385) and (hState = 334)) or
								((vState = 385) and (hState = 335)) or
								((vState = 385) and (hState = 336)) or
								((vState = 385) and (hState = 341)) or
								((vState = 385) and (hState = 357)) or
								((vState = 385) and (hState = 358)) or
								((vState = 385) and (hState = 359)) or
								((vState = 385) and (hState = 385)) or
								((vState = 385) and (hState = 386)) or
								((vState = 385) and (hState = 387)) or
								((vState = 385) and (hState = 392)) or
								((vState = 385) and (hState = 405)) or
								((vState = 385) and (hState = 406)) or
								((vState = 385) and (hState = 428)) or
								((vState = 385) and (hState = 429)) or
								((vState = 385) and (hState = 468)) or
								((vState = 385) and (hState = 469)) or
								((vState = 385) and (hState = 470)) or
								((vState = 385) and (hState = 471)) or
								((vState = 385) and (hState = 472)) or
								((vState = 385) and (hState = 473)) or
								((vState = 385) and (hState = 474)) or
								((vState = 385) and (hState = 490)) or
								((vState = 385) and (hState = 532)) or
								((vState = 385) and (hState = 572)) or
								((vState = 385) and (hState = 583)) or
								((vState = 385) and (hState = 588)) or
								((vState = 386) and (hState = 230)) or
								((vState = 386) and (hState = 231)) or
								((vState = 386) and (hState = 232)) or
								((vState = 386) and (hState = 233)) or
								((vState = 386) and (hState = 234)) or
								((vState = 386) and (hState = 272)) or
								((vState = 386) and (hState = 278)) or
								((vState = 386) and (hState = 279)) or
								((vState = 386) and (hState = 320)) or
								((vState = 386) and (hState = 328)) or
								((vState = 386) and (hState = 329)) or
								((vState = 386) and (hState = 330)) or
								((vState = 386) and (hState = 341)) or
								((vState = 386) and (hState = 359)) or
								((vState = 386) and (hState = 360)) or
								((vState = 386) and (hState = 361)) or
								((vState = 386) and (hState = 362)) or
								((vState = 386) and (hState = 384)) or
								((vState = 386) and (hState = 385)) or
								((vState = 386) and (hState = 392)) or
								((vState = 386) and (hState = 407)) or
								((vState = 386) and (hState = 428)) or
								((vState = 386) and (hState = 429)) or
								((vState = 386) and (hState = 466)) or
								((vState = 386) and (hState = 475)) or
								((vState = 386) and (hState = 476)) or
								((vState = 386) and (hState = 477)) or
								((vState = 386) and (hState = 478)) or
								((vState = 386) and (hState = 479)) or
								((vState = 386) and (hState = 480)) or
								((vState = 386) and (hState = 481)) or
								((vState = 386) and (hState = 482)) or
								((vState = 386) and (hState = 491)) or
								((vState = 386) and (hState = 511)) or
								((vState = 386) and (hState = 532)) or
								((vState = 386) and (hState = 573)) or
								((vState = 386) and (hState = 584)) or
								((vState = 386) and (hState = 588)) or
								((vState = 386) and (hState = 589)) or
								((vState = 387) and (hState = 230)) or
								((vState = 387) and (hState = 231)) or
								((vState = 387) and (hState = 273)) or
								((vState = 387) and (hState = 277)) or
								((vState = 387) and (hState = 320)) or
								((vState = 387) and (hState = 321)) or
								((vState = 387) and (hState = 322)) or
								((vState = 387) and (hState = 323)) or
								((vState = 387) and (hState = 324)) or
								((vState = 387) and (hState = 325)) or
								((vState = 387) and (hState = 330)) or
								((vState = 387) and (hState = 360)) or
								((vState = 387) and (hState = 361)) or
								((vState = 387) and (hState = 362)) or
								((vState = 387) and (hState = 363)) or
								((vState = 387) and (hState = 364)) or
								((vState = 387) and (hState = 379)) or
								((vState = 387) and (hState = 383)) or
								((vState = 387) and (hState = 384)) or
								((vState = 387) and (hState = 392)) or
								((vState = 387) and (hState = 400)) or
								((vState = 387) and (hState = 407)) or
								((vState = 387) and (hState = 428)) or
								((vState = 387) and (hState = 429)) or
								((vState = 387) and (hState = 463)) or
								((vState = 387) and (hState = 464)) or
								((vState = 387) and (hState = 479)) or
								((vState = 387) and (hState = 480)) or
								((vState = 387) and (hState = 481)) or
								((vState = 387) and (hState = 482)) or
								((vState = 387) and (hState = 492)) or
								((vState = 387) and (hState = 512)) or
								((vState = 387) and (hState = 517)) or
								((vState = 387) and (hState = 532)) or
								((vState = 387) and (hState = 574)) or
								((vState = 387) and (hState = 584)) or
								((vState = 387) and (hState = 585)) or
								((vState = 387) and (hState = 586)) or
								((vState = 387) and (hState = 587)) or
								((vState = 387) and (hState = 588)) or
								((vState = 387) and (hState = 589)) or
								((vState = 388) and (hState = 273)) or
								((vState = 388) and (hState = 274)) or
								((vState = 388) and (hState = 320)) or
								((vState = 388) and (hState = 321)) or
								((vState = 388) and (hState = 361)) or
								((vState = 388) and (hState = 362)) or
								((vState = 388) and (hState = 383)) or
								((vState = 388) and (hState = 384)) or
								((vState = 388) and (hState = 392)) or
								((vState = 388) and (hState = 403)) or
								((vState = 388) and (hState = 428)) or
								((vState = 388) and (hState = 458)) or
								((vState = 388) and (hState = 463)) or
								((vState = 388) and (hState = 464)) or
								((vState = 388) and (hState = 479)) or
								((vState = 388) and (hState = 480)) or
								((vState = 388) and (hState = 481)) or
								((vState = 388) and (hState = 482)) or
								((vState = 388) and (hState = 492)) or
								((vState = 388) and (hState = 517)) or
								((vState = 388) and (hState = 532)) or
								((vState = 388) and (hState = 584)) or
								((vState = 388) and (hState = 585)) or
								((vState = 388) and (hState = 586)) or
								((vState = 388) and (hState = 587)) or
								((vState = 388) and (hState = 588)) or
								((vState = 388) and (hState = 589)) or
								((vState = 389) and (hState = 273)) or
								((vState = 389) and (hState = 274)) or
								((vState = 389) and (hState = 275)) or
								((vState = 389) and (hState = 276)) or
								((vState = 389) and (hState = 362)) or
								((vState = 389) and (hState = 383)) or
								((vState = 389) and (hState = 402)) or
								((vState = 389) and (hState = 427)) or
								((vState = 389) and (hState = 428)) or
								((vState = 389) and (hState = 458)) or
								((vState = 389) and (hState = 459)) or
								((vState = 389) and (hState = 460)) or
								((vState = 389) and (hState = 461)) or
								((vState = 389) and (hState = 462)) or
								((vState = 389) and (hState = 463)) or
								((vState = 389) and (hState = 464)) or
								((vState = 389) and (hState = 479)) or
								((vState = 389) and (hState = 480)) or
								((vState = 389) and (hState = 481)) or
								((vState = 389) and (hState = 482)) or
								((vState = 389) and (hState = 492)) or
								((vState = 389) and (hState = 493)) or
								((vState = 389) and (hState = 494)) or
								((vState = 389) and (hState = 495)) or
								((vState = 389) and (hState = 517)) or
								((vState = 389) and (hState = 532)) or
								((vState = 389) and (hState = 569)) or
								((vState = 389) and (hState = 584)) or
								((vState = 389) and (hState = 585)) or
								((vState = 389) and (hState = 586)) or
								((vState = 389) and (hState = 587)) or
								((vState = 389) and (hState = 588)) or
								((vState = 389) and (hState = 589)) or
								((vState = 390) and (hState = 273)) or
								((vState = 390) and (hState = 274)) or
								((vState = 390) and (hState = 275)) or
								((vState = 390) and (hState = 276)) or
								((vState = 390) and (hState = 315)) or
								((vState = 390) and (hState = 316)) or
								((vState = 390) and (hState = 329)) or
								((vState = 390) and (hState = 342)) or
								((vState = 390) and (hState = 362)) or
								((vState = 390) and (hState = 368)) or
								((vState = 390) and (hState = 377)) or
								((vState = 390) and (hState = 381)) or
								((vState = 390) and (hState = 382)) or
								((vState = 390) and (hState = 383)) or
								((vState = 390) and (hState = 402)) or
								((vState = 390) and (hState = 427)) or
								((vState = 390) and (hState = 428)) or
								((vState = 390) and (hState = 457)) or
								((vState = 390) and (hState = 458)) or
								((vState = 390) and (hState = 459)) or
								((vState = 390) and (hState = 460)) or
								((vState = 390) and (hState = 461)) or
								((vState = 390) and (hState = 462)) or
								((vState = 390) and (hState = 463)) or
								((vState = 390) and (hState = 464)) or
								((vState = 390) and (hState = 465)) or
								((vState = 390) and (hState = 466)) or
								((vState = 390) and (hState = 467)) or
								((vState = 390) and (hState = 468)) or
								((vState = 390) and (hState = 469)) or
								((vState = 390) and (hState = 470)) or
								((vState = 390) and (hState = 471)) or
								((vState = 390) and (hState = 472)) or
								((vState = 390) and (hState = 473)) or
								((vState = 390) and (hState = 474)) or
								((vState = 390) and (hState = 475)) or
								((vState = 390) and (hState = 476)) or
								((vState = 390) and (hState = 477)) or
								((vState = 390) and (hState = 478)) or
								((vState = 390) and (hState = 479)) or
								((vState = 390) and (hState = 480)) or
								((vState = 390) and (hState = 481)) or
								((vState = 390) and (hState = 482)) or
								((vState = 390) and (hState = 483)) or
								((vState = 390) and (hState = 484)) or
								((vState = 390) and (hState = 485)) or
								((vState = 390) and (hState = 486)) or
								((vState = 390) and (hState = 487)) or
								((vState = 390) and (hState = 488)) or
								((vState = 390) and (hState = 489)) or
								((vState = 390) and (hState = 490)) or
								((vState = 390) and (hState = 491)) or
								((vState = 390) and (hState = 492)) or
								((vState = 390) and (hState = 493)) or
								((vState = 390) and (hState = 494)) or
								((vState = 390) and (hState = 495)) or
								((vState = 390) and (hState = 496)) or
								((vState = 390) and (hState = 497)) or
								((vState = 390) and (hState = 498)) or
								((vState = 390) and (hState = 499)) or
								((vState = 390) and (hState = 517)) or
								((vState = 390) and (hState = 532)) or
								((vState = 390) and (hState = 569)) or
								((vState = 390) and (hState = 577)) or
								((vState = 390) and (hState = 584)) or
								((vState = 390) and (hState = 585)) or
								((vState = 390) and (hState = 586)) or
								((vState = 390) and (hState = 587)) or
								((vState = 390) and (hState = 588)) or
								((vState = 390) and (hState = 589)) or
								((vState = 391) and (hState = 272)) or
								((vState = 391) and (hState = 277)) or
								((vState = 391) and (hState = 310)) or
								((vState = 391) and (hState = 311)) or
								((vState = 391) and (hState = 312)) or
								((vState = 391) and (hState = 313)) or
								((vState = 391) and (hState = 329)) or
								((vState = 391) and (hState = 340)) or
								((vState = 391) and (hState = 341)) or
								((vState = 391) and (hState = 342)) or
								((vState = 391) and (hState = 343)) or
								((vState = 391) and (hState = 363)) or
								((vState = 391) and (hState = 370)) or
								((vState = 391) and (hState = 371)) or
								((vState = 391) and (hState = 381)) or
								((vState = 391) and (hState = 382)) or
								((vState = 391) and (hState = 383)) or
								((vState = 391) and (hState = 402)) or
								((vState = 391) and (hState = 427)) or
								((vState = 391) and (hState = 428)) or
								((vState = 391) and (hState = 460)) or
								((vState = 391) and (hState = 471)) or
								((vState = 391) and (hState = 491)) or
								((vState = 391) and (hState = 492)) or
								((vState = 391) and (hState = 493)) or
								((vState = 391) and (hState = 494)) or
								((vState = 391) and (hState = 495)) or
								((vState = 391) and (hState = 496)) or
								((vState = 391) and (hState = 497)) or
								((vState = 391) and (hState = 498)) or
								((vState = 391) and (hState = 514)) or
								((vState = 391) and (hState = 515)) or
								((vState = 391) and (hState = 516)) or
								((vState = 391) and (hState = 517)) or
								((vState = 391) and (hState = 532)) or
								((vState = 391) and (hState = 569)) or
								((vState = 391) and (hState = 585)) or
								((vState = 391) and (hState = 586)) or
								((vState = 391) and (hState = 590)) or
								((vState = 392) and (hState = 269)) or
								((vState = 392) and (hState = 278)) or
								((vState = 392) and (hState = 307)) or
								((vState = 392) and (hState = 308)) or
								((vState = 392) and (hState = 329)) or
								((vState = 392) and (hState = 341)) or
								((vState = 392) and (hState = 342)) or
								((vState = 392) and (hState = 343)) or
								((vState = 392) and (hState = 352)) or
								((vState = 392) and (hState = 372)) or
								((vState = 392) and (hState = 381)) or
								((vState = 392) and (hState = 382)) or
								((vState = 392) and (hState = 402)) or
								((vState = 392) and (hState = 403)) or
								((vState = 392) and (hState = 427)) or
								((vState = 392) and (hState = 460)) or
								((vState = 392) and (hState = 491)) or
								((vState = 392) and (hState = 492)) or
								((vState = 392) and (hState = 513)) or
								((vState = 392) and (hState = 514)) or
								((vState = 392) and (hState = 515)) or
								((vState = 392) and (hState = 516)) or
								((vState = 392) and (hState = 517)) or
								((vState = 392) and (hState = 518)) or
								((vState = 392) and (hState = 532)) or
								((vState = 392) and (hState = 542)) or
								((vState = 392) and (hState = 569)) or
								((vState = 392) and (hState = 585)) or
								((vState = 392) and (hState = 586)) or
								((vState = 393) and (hState = 301)) or
								((vState = 393) and (hState = 329)) or
								((vState = 393) and (hState = 342)) or
								((vState = 393) and (hState = 343)) or
								((vState = 393) and (hState = 352)) or
								((vState = 393) and (hState = 380)) or
								((vState = 393) and (hState = 381)) or
								((vState = 393) and (hState = 382)) or
								((vState = 393) and (hState = 427)) or
								((vState = 393) and (hState = 484)) or
								((vState = 393) and (hState = 518)) or
								((vState = 393) and (hState = 532)) or
								((vState = 393) and (hState = 542)) or
								((vState = 393) and (hState = 585)) or
								((vState = 393) and (hState = 586)) or
								((vState = 394) and (hState = 251)) or
								((vState = 394) and (hState = 343)) or
								((vState = 394) and (hState = 344)) or
								((vState = 394) and (hState = 352)) or
								((vState = 394) and (hState = 373)) or
								((vState = 394) and (hState = 374)) or
								((vState = 394) and (hState = 379)) or
								((vState = 394) and (hState = 380)) or
								((vState = 394) and (hState = 401)) or
								((vState = 394) and (hState = 410)) or
								((vState = 394) and (hState = 426)) or
								((vState = 394) and (hState = 427)) or
								((vState = 394) and (hState = 484)) or
								((vState = 394) and (hState = 485)) or
								((vState = 394) and (hState = 486)) or
								((vState = 394) and (hState = 518)) or
								((vState = 394) and (hState = 532)) or
								((vState = 394) and (hState = 542)) or
								((vState = 394) and (hState = 568)) or
								((vState = 394) and (hState = 584)) or
								((vState = 394) and (hState = 585)) or
								((vState = 394) and (hState = 586)) or
								((vState = 395) and (hState = 251)) or
								((vState = 395) and (hState = 343)) or
								((vState = 395) and (hState = 344)) or
								((vState = 395) and (hState = 345)) or
								((vState = 395) and (hState = 352)) or
								((vState = 395) and (hState = 367)) or
								((vState = 395) and (hState = 373)) or
								((vState = 395) and (hState = 374)) or
								((vState = 395) and (hState = 375)) or
								((vState = 395) and (hState = 376)) or
								((vState = 395) and (hState = 377)) or
								((vState = 395) and (hState = 378)) or
								((vState = 395) and (hState = 379)) or
								((vState = 395) and (hState = 380)) or
								((vState = 395) and (hState = 401)) or
								((vState = 395) and (hState = 406)) or
								((vState = 395) and (hState = 410)) or
								((vState = 395) and (hState = 411)) or
								((vState = 395) and (hState = 426)) or
								((vState = 395) and (hState = 427)) or
								((vState = 395) and (hState = 465)) or
								((vState = 395) and (hState = 474)) or
								((vState = 395) and (hState = 484)) or
								((vState = 395) and (hState = 485)) or
								((vState = 395) and (hState = 486)) or
								((vState = 395) and (hState = 501)) or
								((vState = 395) and (hState = 502)) or
								((vState = 395) and (hState = 503)) or
								((vState = 395) and (hState = 504)) or
								((vState = 395) and (hState = 518)) or
								((vState = 395) and (hState = 519)) or
								((vState = 395) and (hState = 542)) or
								((vState = 395) and (hState = 553)) or
								((vState = 395) and (hState = 554)) or
								((vState = 395) and (hState = 568)) or
								((vState = 395) and (hState = 582)) or
								((vState = 395) and (hState = 583)) or
								((vState = 395) and (hState = 584)) or
								((vState = 395) and (hState = 585)) or
								((vState = 395) and (hState = 586)) or
								((vState = 395) and (hState = 594)) or
								((vState = 396) and (hState = 251)) or
								((vState = 396) and (hState = 281)) or
								((vState = 396) and (hState = 299)) or
								((vState = 396) and (hState = 300)) or
								((vState = 396) and (hState = 325)) or
								((vState = 396) and (hState = 326)) or
								((vState = 396) and (hState = 327)) or
								((vState = 396) and (hState = 344)) or
								((vState = 396) and (hState = 345)) or
								((vState = 396) and (hState = 352)) or
								((vState = 396) and (hState = 368)) or
								((vState = 396) and (hState = 372)) or
								((vState = 396) and (hState = 377)) or
								((vState = 396) and (hState = 378)) or
								((vState = 396) and (hState = 379)) or
								((vState = 396) and (hState = 380)) or
								((vState = 396) and (hState = 401)) or
								((vState = 396) and (hState = 410)) or
								((vState = 396) and (hState = 411)) or
								((vState = 396) and (hState = 412)) or
								((vState = 396) and (hState = 413)) or
								((vState = 396) and (hState = 414)) or
								((vState = 396) and (hState = 415)) or
								((vState = 396) and (hState = 416)) or
								((vState = 396) and (hState = 417)) or
								((vState = 396) and (hState = 418)) or
								((vState = 396) and (hState = 419)) or
								((vState = 396) and (hState = 420)) or
								((vState = 396) and (hState = 421)) or
								((vState = 396) and (hState = 422)) or
								((vState = 396) and (hState = 423)) or
								((vState = 396) and (hState = 424)) or
								((vState = 396) and (hState = 425)) or
								((vState = 396) and (hState = 426)) or
								((vState = 396) and (hState = 427)) or
								((vState = 396) and (hState = 428)) or
								((vState = 396) and (hState = 429)) or
								((vState = 396) and (hState = 430)) or
								((vState = 396) and (hState = 431)) or
								((vState = 396) and (hState = 432)) or
								((vState = 396) and (hState = 433)) or
								((vState = 396) and (hState = 434)) or
								((vState = 396) and (hState = 435)) or
								((vState = 396) and (hState = 436)) or
								((vState = 396) and (hState = 437)) or
								((vState = 396) and (hState = 438)) or
								((vState = 396) and (hState = 463)) or
								((vState = 396) and (hState = 464)) or
								((vState = 396) and (hState = 475)) or
								((vState = 396) and (hState = 480)) or
								((vState = 396) and (hState = 481)) or
								((vState = 396) and (hState = 486)) or
								((vState = 396) and (hState = 495)) or
								((vState = 396) and (hState = 496)) or
								((vState = 396) and (hState = 497)) or
								((vState = 396) and (hState = 498)) or
								((vState = 396) and (hState = 503)) or
								((vState = 396) and (hState = 504)) or
								((vState = 396) and (hState = 518)) or
								((vState = 396) and (hState = 519)) or
								((vState = 396) and (hState = 531)) or
								((vState = 396) and (hState = 542)) or
								((vState = 396) and (hState = 553)) or
								((vState = 396) and (hState = 554)) or
								((vState = 396) and (hState = 568)) or
								((vState = 396) and (hState = 582)) or
								((vState = 396) and (hState = 583)) or
								((vState = 396) and (hState = 595)) or
								((vState = 397) and (hState = 251)) or
								((vState = 397) and (hState = 282)) or
								((vState = 397) and (hState = 299)) or
								((vState = 397) and (hState = 300)) or
								((vState = 397) and (hState = 325)) or
								((vState = 397) and (hState = 326)) or
								((vState = 397) and (hState = 327)) or
								((vState = 397) and (hState = 345)) or
								((vState = 397) and (hState = 346)) or
								((vState = 397) and (hState = 370)) or
								((vState = 397) and (hState = 371)) or
								((vState = 397) and (hState = 377)) or
								((vState = 397) and (hState = 400)) or
								((vState = 397) and (hState = 412)) or
								((vState = 397) and (hState = 425)) or
								((vState = 397) and (hState = 443)) or
								((vState = 397) and (hState = 444)) or
								((vState = 397) and (hState = 463)) or
								((vState = 397) and (hState = 464)) or
								((vState = 397) and (hState = 475)) or
								((vState = 397) and (hState = 476)) or
								((vState = 397) and (hState = 477)) or
								((vState = 397) and (hState = 478)) or
								((vState = 397) and (hState = 486)) or
								((vState = 397) and (hState = 487)) or
								((vState = 397) and (hState = 488)) or
								((vState = 397) and (hState = 489)) or
								((vState = 397) and (hState = 490)) or
								((vState = 397) and (hState = 491)) or
								((vState = 397) and (hState = 492)) or
								((vState = 397) and (hState = 518)) or
								((vState = 397) and (hState = 519)) or
								((vState = 397) and (hState = 520)) or
								((vState = 397) and (hState = 531)) or
								((vState = 397) and (hState = 542)) or
								((vState = 397) and (hState = 553)) or
								((vState = 397) and (hState = 554)) or
								((vState = 397) and (hState = 582)) or
								((vState = 397) and (hState = 583)) or
								((vState = 398) and (hState = 251)) or
								((vState = 398) and (hState = 299)) or
								((vState = 398) and (hState = 300)) or
								((vState = 398) and (hState = 326)) or
								((vState = 398) and (hState = 327)) or
								((vState = 398) and (hState = 345)) or
								((vState = 398) and (hState = 346)) or
								((vState = 398) and (hState = 370)) or
								((vState = 398) and (hState = 371)) or
								((vState = 398) and (hState = 381)) or
								((vState = 398) and (hState = 400)) or
								((vState = 398) and (hState = 412)) or
								((vState = 398) and (hState = 425)) or
								((vState = 398) and (hState = 474)) or
								((vState = 398) and (hState = 475)) or
								((vState = 398) and (hState = 476)) or
								((vState = 398) and (hState = 477)) or
								((vState = 398) and (hState = 478)) or
								((vState = 398) and (hState = 485)) or
								((vState = 398) and (hState = 486)) or
								((vState = 398) and (hState = 487)) or
								((vState = 398) and (hState = 488)) or
								((vState = 398) and (hState = 518)) or
								((vState = 398) and (hState = 531)) or
								((vState = 398) and (hState = 538)) or
								((vState = 398) and (hState = 553)) or
								((vState = 398) and (hState = 554)) or
								((vState = 398) and (hState = 586)) or
								((vState = 399) and (hState = 252)) or
								((vState = 399) and (hState = 299)) or
								((vState = 399) and (hState = 300)) or
								((vState = 399) and (hState = 326)) or
								((vState = 399) and (hState = 346)) or
								((vState = 399) and (hState = 351)) or
								((vState = 399) and (hState = 370)) or
								((vState = 399) and (hState = 371)) or
								((vState = 399) and (hState = 400)) or
								((vState = 399) and (hState = 412)) or
								((vState = 399) and (hState = 425)) or
								((vState = 399) and (hState = 474)) or
								((vState = 399) and (hState = 475)) or
								((vState = 399) and (hState = 476)) or
								((vState = 399) and (hState = 477)) or
								((vState = 399) and (hState = 478)) or
								((vState = 399) and (hState = 479)) or
								((vState = 399) and (hState = 522)) or
								((vState = 399) and (hState = 531)) or
								((vState = 399) and (hState = 537)) or
								((vState = 399) and (hState = 553)) or
								((vState = 399) and (hState = 567)) or
								((vState = 399) and (hState = 585)) or
								((vState = 399) and (hState = 586)) or
								((vState = 400) and (hState = 299)) or
								((vState = 400) and (hState = 300)) or
								((vState = 400) and (hState = 326)) or
								((vState = 400) and (hState = 351)) or
								((vState = 400) and (hState = 425)) or
								((vState = 400) and (hState = 461)) or
								((vState = 400) and (hState = 465)) or
								((vState = 400) and (hState = 470)) or
								((vState = 400) and (hState = 471)) or
								((vState = 400) and (hState = 472)) or
								((vState = 400) and (hState = 473)) or
								((vState = 400) and (hState = 474)) or
								((vState = 400) and (hState = 475)) or
								((vState = 400) and (hState = 478)) or
								((vState = 400) and (hState = 479)) or
								((vState = 400) and (hState = 480)) or
								((vState = 400) and (hState = 522)) or
								((vState = 400) and (hState = 523)) or
								((vState = 400) and (hState = 531)) or
								((vState = 400) and (hState = 532)) or
								((vState = 400) and (hState = 537)) or
								((vState = 400) and (hState = 552)) or
								((vState = 400) and (hState = 553)) or
								((vState = 400) and (hState = 567)) or
								((vState = 400) and (hState = 586)) or
								((vState = 401) and (hState = 299)) or
								((vState = 401) and (hState = 300)) or
								((vState = 401) and (hState = 326)) or
								((vState = 401) and (hState = 347)) or
								((vState = 401) and (hState = 351)) or
								((vState = 401) and (hState = 368)) or
								((vState = 401) and (hState = 373)) or
								((vState = 401) and (hState = 374)) or
								((vState = 401) and (hState = 385)) or
								((vState = 401) and (hState = 386)) or
								((vState = 401) and (hState = 387)) or
								((vState = 401) and (hState = 413)) or
								((vState = 401) and (hState = 458)) or
								((vState = 401) and (hState = 459)) or
								((vState = 401) and (hState = 460)) or
								((vState = 401) and (hState = 461)) or
								((vState = 401) and (hState = 465)) or
								((vState = 401) and (hState = 466)) or
								((vState = 401) and (hState = 467)) or
								((vState = 401) and (hState = 468)) or
								((vState = 401) and (hState = 469)) or
								((vState = 401) and (hState = 470)) or
								((vState = 401) and (hState = 471)) or
								((vState = 401) and (hState = 472)) or
								((vState = 401) and (hState = 473)) or
								((vState = 401) and (hState = 474)) or
								((vState = 401) and (hState = 475)) or
								((vState = 401) and (hState = 479)) or
								((vState = 401) and (hState = 480)) or
								((vState = 401) and (hState = 490)) or
								((vState = 401) and (hState = 523)) or
								((vState = 401) and (hState = 524)) or
								((vState = 401) and (hState = 531)) or
								((vState = 401) and (hState = 532)) or
								((vState = 401) and (hState = 533)) or
								((vState = 401) and (hState = 534)) or
								((vState = 401) and (hState = 537)) or
								((vState = 401) and (hState = 541)) or
								((vState = 401) and (hState = 552)) or
								((vState = 401) and (hState = 553)) or
								((vState = 401) and (hState = 567)) or
								((vState = 401) and (hState = 578)) or
								((vState = 402) and (hState = 298)) or
								((vState = 402) and (hState = 299)) or
								((vState = 402) and (hState = 300)) or
								((vState = 402) and (hState = 326)) or
								((vState = 402) and (hState = 327)) or
								((vState = 402) and (hState = 347)) or
								((vState = 402) and (hState = 351)) or
								((vState = 402) and (hState = 373)) or
								((vState = 402) and (hState = 374)) or
								((vState = 402) and (hState = 379)) or
								((vState = 402) and (hState = 388)) or
								((vState = 402) and (hState = 413)) or
								((vState = 402) and (hState = 458)) or
								((vState = 402) and (hState = 459)) or
								((vState = 402) and (hState = 460)) or
								((vState = 402) and (hState = 461)) or
								((vState = 402) and (hState = 462)) or
								((vState = 402) and (hState = 463)) or
								((vState = 402) and (hState = 464)) or
								((vState = 402) and (hState = 465)) or
								((vState = 402) and (hState = 466)) or
								((vState = 402) and (hState = 467)) or
								((vState = 402) and (hState = 468)) or
								((vState = 402) and (hState = 469)) or
								((vState = 402) and (hState = 480)) or
								((vState = 402) and (hState = 511)) or
								((vState = 402) and (hState = 519)) or
								((vState = 402) and (hState = 524)) or
								((vState = 402) and (hState = 525)) or
								((vState = 402) and (hState = 531)) or
								((vState = 402) and (hState = 532)) or
								((vState = 402) and (hState = 541)) or
								((vState = 402) and (hState = 552)) or
								((vState = 402) and (hState = 553)) or
								((vState = 402) and (hState = 567)) or
								((vState = 402) and (hState = 587)) or
								((vState = 402) and (hState = 588)) or
								((vState = 403) and (hState = 287)) or
								((vState = 403) and (hState = 298)) or
								((vState = 403) and (hState = 299)) or
								((vState = 403) and (hState = 300)) or
								((vState = 403) and (hState = 326)) or
								((vState = 403) and (hState = 327)) or
								((vState = 403) and (hState = 350)) or
								((vState = 403) and (hState = 367)) or
								((vState = 403) and (hState = 379)) or
								((vState = 403) and (hState = 395)) or
								((vState = 403) and (hState = 424)) or
								((vState = 403) and (hState = 458)) or
								((vState = 403) and (hState = 459)) or
								((vState = 403) and (hState = 460)) or
								((vState = 403) and (hState = 461)) or
								((vState = 403) and (hState = 462)) or
								((vState = 403) and (hState = 468)) or
								((vState = 403) and (hState = 469)) or
								((vState = 403) and (hState = 491)) or
								((vState = 403) and (hState = 512)) or
								((vState = 403) and (hState = 519)) or
								((vState = 403) and (hState = 524)) or
								((vState = 403) and (hState = 525)) or
								((vState = 403) and (hState = 526)) or
								((vState = 403) and (hState = 531)) or
								((vState = 403) and (hState = 536)) or
								((vState = 403) and (hState = 541)) or
								((vState = 403) and (hState = 552)) or
								((vState = 403) and (hState = 553)) or
								((vState = 403) and (hState = 577)) or
								((vState = 403) and (hState = 587)) or
								((vState = 403) and (hState = 588)) or
								((vState = 403) and (hState = 589)) or
								((vState = 404) and (hState = 298)) or
								((vState = 404) and (hState = 299)) or
								((vState = 404) and (hState = 300)) or
								((vState = 404) and (hState = 350)) or
								((vState = 404) and (hState = 366)) or
								((vState = 404) and (hState = 379)) or
								((vState = 404) and (hState = 395)) or
								((vState = 404) and (hState = 423)) or
								((vState = 404) and (hState = 458)) or
								((vState = 404) and (hState = 469)) or
								((vState = 404) and (hState = 491)) or
								((vState = 404) and (hState = 519)) or
								((vState = 404) and (hState = 525)) or
								((vState = 404) and (hState = 526)) or
								((vState = 404) and (hState = 527)) or
								((vState = 404) and (hState = 531)) or
								((vState = 404) and (hState = 541)) or
								((vState = 404) and (hState = 552)) or
								((vState = 404) and (hState = 553)) or
								((vState = 404) and (hState = 587)) or
								((vState = 404) and (hState = 588)) or
								((vState = 404) and (hState = 589)) or
								((vState = 405) and (hState = 300)) or
								((vState = 405) and (hState = 329)) or
								((vState = 405) and (hState = 350)) or
								((vState = 405) and (hState = 371)) or
								((vState = 405) and (hState = 379)) or
								((vState = 405) and (hState = 394)) or
								((vState = 405) and (hState = 395)) or
								((vState = 405) and (hState = 396)) or
								((vState = 405) and (hState = 397)) or
								((vState = 405) and (hState = 423)) or
								((vState = 405) and (hState = 470)) or
								((vState = 405) and (hState = 481)) or
								((vState = 405) and (hState = 492)) or
								((vState = 405) and (hState = 493)) or
								((vState = 405) and (hState = 519)) or
								((vState = 405) and (hState = 525)) or
								((vState = 405) and (hState = 526)) or
								((vState = 405) and (hState = 527)) or
								((vState = 405) and (hState = 528)) or
								((vState = 405) and (hState = 529)) or
								((vState = 405) and (hState = 530)) or
								((vState = 405) and (hState = 541)) or
								((vState = 405) and (hState = 551)) or
								((vState = 405) and (hState = 552)) or
								((vState = 405) and (hState = 553)) or
								((vState = 405) and (hState = 587)) or
								((vState = 405) and (hState = 588)) or
								((vState = 405) and (hState = 589)) or
								((vState = 405) and (hState = 590)) or
								((vState = 406) and (hState = 325)) or
								((vState = 406) and (hState = 329)) or
								((vState = 406) and (hState = 350)) or
								((vState = 406) and (hState = 371)) or
								((vState = 406) and (hState = 377)) or
								((vState = 406) and (hState = 378)) or
								((vState = 406) and (hState = 379)) or
								((vState = 406) and (hState = 394)) or
								((vState = 406) and (hState = 395)) or
								((vState = 406) and (hState = 396)) or
								((vState = 406) and (hState = 397)) or
								((vState = 406) and (hState = 423)) or
								((vState = 406) and (hState = 470)) or
								((vState = 406) and (hState = 475)) or
								((vState = 406) and (hState = 476)) or
								((vState = 406) and (hState = 477)) or
								((vState = 406) and (hState = 478)) or
								((vState = 406) and (hState = 479)) or
								((vState = 406) and (hState = 480)) or
								((vState = 406) and (hState = 481)) or
								((vState = 406) and (hState = 482)) or
								((vState = 406) and (hState = 483)) or
								((vState = 406) and (hState = 484)) or
								((vState = 406) and (hState = 485)) or
								((vState = 406) and (hState = 486)) or
								((vState = 406) and (hState = 487)) or
								((vState = 406) and (hState = 488)) or
								((vState = 406) and (hState = 492)) or
								((vState = 406) and (hState = 493)) or
								((vState = 406) and (hState = 502)) or
								((vState = 406) and (hState = 503)) or
								((vState = 406) and (hState = 519)) or
								((vState = 406) and (hState = 525)) or
								((vState = 406) and (hState = 526)) or
								((vState = 406) and (hState = 527)) or
								((vState = 406) and (hState = 528)) or
								((vState = 406) and (hState = 529)) or
								((vState = 406) and (hState = 530)) or
								((vState = 406) and (hState = 535)) or
								((vState = 406) and (hState = 541)) or
								((vState = 406) and (hState = 550)) or
								((vState = 406) and (hState = 551)) or
								((vState = 406) and (hState = 552)) or
								((vState = 406) and (hState = 553)) or
								((vState = 406) and (hState = 574)) or
								((vState = 406) and (hState = 587)) or
								((vState = 406) and (hState = 588)) or
								((vState = 406) and (hState = 589)) or
								((vState = 406) and (hState = 590)) or
								((vState = 406) and (hState = 591)) or
								((vState = 407) and (hState = 256)) or
								((vState = 407) and (hState = 297)) or
								((vState = 407) and (hState = 325)) or
								((vState = 407) and (hState = 350)) or
								((vState = 407) and (hState = 378)) or
								((vState = 407) and (hState = 379)) or
								((vState = 407) and (hState = 395)) or
								((vState = 407) and (hState = 396)) or
								((vState = 407) and (hState = 397)) or
								((vState = 407) and (hState = 416)) or
								((vState = 407) and (hState = 423)) or
								((vState = 407) and (hState = 455)) or
								((vState = 407) and (hState = 470)) or
								((vState = 407) and (hState = 475)) or
								((vState = 407) and (hState = 476)) or
								((vState = 407) and (hState = 477)) or
								((vState = 407) and (hState = 478)) or
								((vState = 407) and (hState = 479)) or
								((vState = 407) and (hState = 480)) or
								((vState = 407) and (hState = 481)) or
								((vState = 407) and (hState = 482)) or
								((vState = 407) and (hState = 483)) or
								((vState = 407) and (hState = 484)) or
								((vState = 407) and (hState = 485)) or
								((vState = 407) and (hState = 506)) or
								((vState = 407) and (hState = 517)) or
								((vState = 407) and (hState = 518)) or
								((vState = 407) and (hState = 519)) or
								((vState = 407) and (hState = 525)) or
								((vState = 407) and (hState = 526)) or
								((vState = 407) and (hState = 527)) or
								((vState = 407) and (hState = 530)) or
								((vState = 407) and (hState = 547)) or
								((vState = 407) and (hState = 551)) or
								((vState = 407) and (hState = 552)) or
								((vState = 407) and (hState = 553)) or
								((vState = 407) and (hState = 573)) or
								((vState = 407) and (hState = 587)) or
								((vState = 407) and (hState = 588)) or
								((vState = 407) and (hState = 589)) or
								((vState = 407) and (hState = 593)) or
								((vState = 408) and (hState = 257)) or
								((vState = 408) and (hState = 297)) or
								((vState = 408) and (hState = 298)) or
								((vState = 408) and (hState = 299)) or
								((vState = 408) and (hState = 325)) or
								((vState = 408) and (hState = 330)) or
								((vState = 408) and (hState = 350)) or
								((vState = 408) and (hState = 363)) or
								((vState = 408) and (hState = 379)) or
								((vState = 408) and (hState = 395)) or
								((vState = 408) and (hState = 396)) or
								((vState = 408) and (hState = 416)) or
								((vState = 408) and (hState = 422)) or
								((vState = 408) and (hState = 423)) or
								((vState = 408) and (hState = 454)) or
								((vState = 408) and (hState = 466)) or
								((vState = 408) and (hState = 467)) or
								((vState = 408) and (hState = 468)) or
								((vState = 408) and (hState = 469)) or
								((vState = 408) and (hState = 470)) or
								((vState = 408) and (hState = 471)) or
								((vState = 408) and (hState = 485)) or
								((vState = 408) and (hState = 508)) or
								((vState = 408) and (hState = 517)) or
								((vState = 408) and (hState = 525)) or
								((vState = 408) and (hState = 526)) or
								((vState = 408) and (hState = 527)) or
								((vState = 408) and (hState = 530)) or
								((vState = 408) and (hState = 531)) or
								((vState = 408) and (hState = 532)) or
								((vState = 408) and (hState = 533)) or
								((vState = 408) and (hState = 540)) or
								((vState = 408) and (hState = 546)) or
								((vState = 408) and (hState = 551)) or
								((vState = 408) and (hState = 552)) or
								((vState = 408) and (hState = 553)) or
								((vState = 408) and (hState = 587)) or
								((vState = 408) and (hState = 588)) or
								((vState = 408) and (hState = 589)) or
								((vState = 408) and (hState = 594)) or
								((vState = 409) and (hState = 257)) or
								((vState = 409) and (hState = 297)) or
								((vState = 409) and (hState = 298)) or
								((vState = 409) and (hState = 299)) or
								((vState = 409) and (hState = 325)) or
								((vState = 409) and (hState = 330)) or
								((vState = 409) and (hState = 379)) or
								((vState = 409) and (hState = 395)) or
								((vState = 409) and (hState = 422)) or
								((vState = 409) and (hState = 454)) or
								((vState = 409) and (hState = 470)) or
								((vState = 409) and (hState = 485)) or
								((vState = 409) and (hState = 530)) or
								((vState = 409) and (hState = 531)) or
								((vState = 409) and (hState = 532)) or
								((vState = 409) and (hState = 533)) or
								((vState = 409) and (hState = 540)) or
								((vState = 409) and (hState = 551)) or
								((vState = 409) and (hState = 552)) or
								((vState = 409) and (hState = 587)) or
								((vState = 409) and (hState = 588)) or
								((vState = 409) and (hState = 589)) or
								((vState = 410) and (hState = 297)) or
								((vState = 410) and (hState = 298)) or
								((vState = 410) and (hState = 299)) or
								((vState = 410) and (hState = 362)) or
								((vState = 410) and (hState = 379)) or
								((vState = 410) and (hState = 380)) or
								((vState = 410) and (hState = 381)) or
								((vState = 410) and (hState = 395)) or
								((vState = 410) and (hState = 422)) or
								((vState = 410) and (hState = 453)) or
								((vState = 410) and (hState = 454)) or
								((vState = 410) and (hState = 470)) or
								((vState = 410) and (hState = 485)) or
								((vState = 410) and (hState = 511)) or
								((vState = 410) and (hState = 514)) or
								((vState = 410) and (hState = 521)) or
								((vState = 410) and (hState = 522)) or
								((vState = 410) and (hState = 529)) or
								((vState = 410) and (hState = 530)) or
								((vState = 410) and (hState = 540)) or
								((vState = 410) and (hState = 550)) or
								((vState = 410) and (hState = 551)) or
								((vState = 410) and (hState = 552)) or
								((vState = 411) and (hState = 292)) or
								((vState = 411) and (hState = 297)) or
								((vState = 411) and (hState = 298)) or
								((vState = 411) and (hState = 299)) or
								((vState = 411) and (hState = 312)) or
								((vState = 411) and (hState = 313)) or
								((vState = 411) and (hState = 324)) or
								((vState = 411) and (hState = 331)) or
								((vState = 411) and (hState = 362)) or
								((vState = 411) and (hState = 379)) or
								((vState = 411) and (hState = 380)) or
								((vState = 411) and (hState = 381)) or
								((vState = 411) and (hState = 382)) or
								((vState = 411) and (hState = 395)) or
								((vState = 411) and (hState = 417)) or
								((vState = 411) and (hState = 422)) or
								((vState = 411) and (hState = 449)) or
								((vState = 411) and (hState = 450)) or
								((vState = 411) and (hState = 451)) or
								((vState = 411) and (hState = 452)) or
								((vState = 411) and (hState = 453)) or
								((vState = 411) and (hState = 454)) or
								((vState = 411) and (hState = 470)) or
								((vState = 411) and (hState = 485)) or
								((vState = 411) and (hState = 486)) or
								((vState = 411) and (hState = 496)) or
								((vState = 411) and (hState = 511)) or
								((vState = 411) and (hState = 512)) or
								((vState = 411) and (hState = 513)) or
								((vState = 411) and (hState = 514)) or
								((vState = 411) and (hState = 521)) or
								((vState = 411) and (hState = 522)) or
								((vState = 411) and (hState = 529)) or
								((vState = 411) and (hState = 530)) or
								((vState = 411) and (hState = 540)) or
								((vState = 411) and (hState = 550)) or
								((vState = 411) and (hState = 551)) or
								((vState = 411) and (hState = 552)) or
								((vState = 411) and (hState = 563)) or
								((vState = 412) and (hState = 293)) or
								((vState = 412) and (hState = 294)) or
								((vState = 412) and (hState = 295)) or
								((vState = 412) and (hState = 296)) or
								((vState = 412) and (hState = 297)) or
								((vState = 412) and (hState = 298)) or
								((vState = 412) and (hState = 299)) or
								((vState = 412) and (hState = 312)) or
								((vState = 412) and (hState = 313)) or
								((vState = 412) and (hState = 324)) or
								((vState = 412) and (hState = 331)) or
								((vState = 412) and (hState = 365)) or
								((vState = 412) and (hState = 366)) or
								((vState = 412) and (hState = 367)) or
								((vState = 412) and (hState = 381)) or
								((vState = 412) and (hState = 382)) or
								((vState = 412) and (hState = 383)) or
								((vState = 412) and (hState = 395)) or
								((vState = 412) and (hState = 417)) or
								((vState = 412) and (hState = 422)) or
								((vState = 412) and (hState = 441)) or
								((vState = 412) and (hState = 442)) or
								((vState = 412) and (hState = 443)) or
								((vState = 412) and (hState = 444)) or
								((vState = 412) and (hState = 445)) or
								((vState = 412) and (hState = 450)) or
								((vState = 412) and (hState = 451)) or
								((vState = 412) and (hState = 470)) or
								((vState = 412) and (hState = 485)) or
								((vState = 412) and (hState = 486)) or
								((vState = 412) and (hState = 487)) or
								((vState = 412) and (hState = 511)) or
								((vState = 412) and (hState = 516)) or
								((vState = 412) and (hState = 517)) or
								((vState = 412) and (hState = 520)) or
								((vState = 412) and (hState = 529)) or
								((vState = 412) and (hState = 530)) or
								((vState = 412) and (hState = 540)) or
								((vState = 412) and (hState = 541)) or
								((vState = 412) and (hState = 542)) or
								((vState = 412) and (hState = 550)) or
								((vState = 412) and (hState = 551)) or
								((vState = 412) and (hState = 552)) or
								((vState = 412) and (hState = 563)) or
								((vState = 412) and (hState = 569)) or
								((vState = 412) and (hState = 590)) or
								((vState = 413) and (hState = 260)) or
								((vState = 413) and (hState = 294)) or
								((vState = 413) and (hState = 295)) or
								((vState = 413) and (hState = 299)) or
								((vState = 413) and (hState = 312)) or
								((vState = 413) and (hState = 313)) or
								((vState = 413) and (hState = 314)) or
								((vState = 413) and (hState = 324)) or
								((vState = 413) and (hState = 366)) or
								((vState = 413) and (hState = 367)) or
								((vState = 413) and (hState = 384)) or
								((vState = 413) and (hState = 418)) or
								((vState = 413) and (hState = 419)) or
								((vState = 413) and (hState = 420)) or
								((vState = 413) and (hState = 421)) or
								((vState = 413) and (hState = 438)) or
								((vState = 413) and (hState = 450)) or
								((vState = 413) and (hState = 470)) or
								((vState = 413) and (hState = 485)) or
								((vState = 413) and (hState = 497)) or
								((vState = 413) and (hState = 517)) or
								((vState = 413) and (hState = 518)) or
								((vState = 413) and (hState = 519)) or
								((vState = 413) and (hState = 520)) or
								((vState = 413) and (hState = 530)) or
								((vState = 413) and (hState = 540)) or
								((vState = 413) and (hState = 541)) or
								((vState = 413) and (hState = 550)) or
								((vState = 413) and (hState = 551)) or
								((vState = 413) and (hState = 552)) or
								((vState = 413) and (hState = 562)) or
								((vState = 413) and (hState = 563)) or
								((vState = 413) and (hState = 588)) or
								((vState = 413) and (hState = 589)) or
								((vState = 413) and (hState = 590)) or
								((vState = 413) and (hState = 599)) or
								((vState = 414) and (hState = 294)) or
								((vState = 414) and (hState = 295)) or
								((vState = 414) and (hState = 299)) or
								((vState = 414) and (hState = 366)) or
								((vState = 414) and (hState = 367)) or
								((vState = 414) and (hState = 385)) or
								((vState = 414) and (hState = 396)) or
								((vState = 414) and (hState = 418)) or
								((vState = 414) and (hState = 419)) or
								((vState = 414) and (hState = 420)) or
								((vState = 414) and (hState = 438)) or
								((vState = 414) and (hState = 470)) or
								((vState = 414) and (hState = 485)) or
								((vState = 414) and (hState = 517)) or
								((vState = 414) and (hState = 521)) or
								((vState = 414) and (hState = 530)) or
								((vState = 414) and (hState = 549)) or
								((vState = 414) and (hState = 550)) or
								((vState = 414) and (hState = 551)) or
								((vState = 414) and (hState = 552)) or
								((vState = 414) and (hState = 562)) or
								((vState = 414) and (hState = 563)) or
								((vState = 414) and (hState = 588)) or
								((vState = 414) and (hState = 589)) or
								((vState = 414) and (hState = 590)) or
								((vState = 415) and (hState = 294)) or
								((vState = 415) and (hState = 295)) or
								((vState = 415) and (hState = 296)) or
								((vState = 415) and (hState = 299)) or
								((vState = 415) and (hState = 386)) or
								((vState = 415) and (hState = 396)) or
								((vState = 415) and (hState = 420)) or
								((vState = 415) and (hState = 438)) or
								((vState = 415) and (hState = 485)) or
								((vState = 415) and (hState = 506)) or
								((vState = 415) and (hState = 521)) or
								((vState = 415) and (hState = 522)) or
								((vState = 415) and (hState = 530)) or
								((vState = 415) and (hState = 549)) or
								((vState = 415) and (hState = 550)) or
								((vState = 415) and (hState = 551)) or
								((vState = 415) and (hState = 552)) or
								((vState = 415) and (hState = 562)) or
								((vState = 415) and (hState = 588)) or
								((vState = 416) and (hState = 261)) or
								((vState = 416) and (hState = 294)) or
								((vState = 416) and (hState = 295)) or
								((vState = 416) and (hState = 296)) or
								((vState = 416) and (hState = 297)) or
								((vState = 416) and (hState = 298)) or
								((vState = 416) and (hState = 299)) or
								((vState = 416) and (hState = 315)) or
								((vState = 416) and (hState = 333)) or
								((vState = 416) and (hState = 341)) or
								((vState = 416) and (hState = 342)) or
								((vState = 416) and (hState = 343)) or
								((vState = 416) and (hState = 344)) or
								((vState = 416) and (hState = 364)) or
								((vState = 416) and (hState = 386)) or
								((vState = 416) and (hState = 387)) or
								((vState = 416) and (hState = 396)) or
								((vState = 416) and (hState = 420)) or
								((vState = 416) and (hState = 438)) or
								((vState = 416) and (hState = 448)) or
								((vState = 416) and (hState = 485)) or
								((vState = 416) and (hState = 490)) or
								((vState = 416) and (hState = 505)) or
								((vState = 416) and (hState = 506)) or
								((vState = 416) and (hState = 515)) or
								((vState = 416) and (hState = 522)) or
								((vState = 416) and (hState = 523)) or
								((vState = 416) and (hState = 524)) or
								((vState = 416) and (hState = 530)) or
								((vState = 416) and (hState = 531)) or
								((vState = 416) and (hState = 537)) or
								((vState = 416) and (hState = 538)) or
								((vState = 416) and (hState = 549)) or
								((vState = 416) and (hState = 550)) or
								((vState = 416) and (hState = 551)) or
								((vState = 416) and (hState = 552)) or
								((vState = 416) and (hState = 562)) or
								((vState = 416) and (hState = 567)) or
								((vState = 416) and (hState = 588)) or
								((vState = 417) and (hState = 293)) or
								((vState = 417) and (hState = 294)) or
								((vState = 417) and (hState = 295)) or
								((vState = 417) and (hState = 296)) or
								((vState = 417) and (hState = 297)) or
								((vState = 417) and (hState = 298)) or
								((vState = 417) and (hState = 299)) or
								((vState = 417) and (hState = 310)) or
								((vState = 417) and (hState = 334)) or
								((vState = 417) and (hState = 338)) or
								((vState = 417) and (hState = 345)) or
								((vState = 417) and (hState = 346)) or
								((vState = 417) and (hState = 347)) or
								((vState = 417) and (hState = 363)) or
								((vState = 417) and (hState = 371)) or
								((vState = 417) and (hState = 388)) or
								((vState = 417) and (hState = 396)) or
								((vState = 417) and (hState = 420)) or
								((vState = 417) and (hState = 438)) or
								((vState = 417) and (hState = 448)) or
								((vState = 417) and (hState = 469)) or
								((vState = 417) and (hState = 485)) or
								((vState = 417) and (hState = 491)) or
								((vState = 417) and (hState = 514)) or
								((vState = 417) and (hState = 522)) or
								((vState = 417) and (hState = 527)) or
								((vState = 417) and (hState = 530)) or
								((vState = 417) and (hState = 531)) or
								((vState = 417) and (hState = 536)) or
								((vState = 417) and (hState = 537)) or
								((vState = 417) and (hState = 538)) or
								((vState = 417) and (hState = 548)) or
								((vState = 417) and (hState = 549)) or
								((vState = 417) and (hState = 550)) or
								((vState = 417) and (hState = 551)) or
								((vState = 417) and (hState = 552)) or
								((vState = 417) and (hState = 561)) or
								((vState = 417) and (hState = 562)) or
								((vState = 417) and (hState = 567)) or
								((vState = 417) and (hState = 588)) or
								((vState = 418) and (hState = 262)) or
								((vState = 418) and (hState = 292)) or
								((vState = 418) and (hState = 293)) or
								((vState = 418) and (hState = 294)) or
								((vState = 418) and (hState = 295)) or
								((vState = 418) and (hState = 296)) or
								((vState = 418) and (hState = 297)) or
								((vState = 418) and (hState = 298)) or
								((vState = 418) and (hState = 299)) or
								((vState = 418) and (hState = 310)) or
								((vState = 418) and (hState = 334)) or
								((vState = 418) and (hState = 335)) or
								((vState = 418) and (hState = 345)) or
								((vState = 418) and (hState = 346)) or
								((vState = 418) and (hState = 347)) or
								((vState = 418) and (hState = 373)) or
								((vState = 418) and (hState = 382)) or
								((vState = 418) and (hState = 389)) or
								((vState = 418) and (hState = 396)) or
								((vState = 418) and (hState = 420)) or
								((vState = 418) and (hState = 438)) or
								((vState = 418) and (hState = 447)) or
								((vState = 418) and (hState = 448)) or
								((vState = 418) and (hState = 449)) or
								((vState = 418) and (hState = 450)) or
								((vState = 418) and (hState = 451)) or
								((vState = 418) and (hState = 452)) or
								((vState = 418) and (hState = 453)) or
								((vState = 418) and (hState = 454)) or
								((vState = 418) and (hState = 455)) or
								((vState = 418) and (hState = 456)) or
								((vState = 418) and (hState = 469)) or
								((vState = 418) and (hState = 485)) or
								((vState = 418) and (hState = 492)) or
								((vState = 418) and (hState = 501)) or
								((vState = 418) and (hState = 502)) or
								((vState = 418) and (hState = 522)) or
								((vState = 418) and (hState = 529)) or
								((vState = 418) and (hState = 530)) or
								((vState = 418) and (hState = 531)) or
								((vState = 418) and (hState = 532)) or
								((vState = 418) and (hState = 533)) or
								((vState = 418) and (hState = 534)) or
								((vState = 418) and (hState = 535)) or
								((vState = 418) and (hState = 547)) or
								((vState = 418) and (hState = 548)) or
								((vState = 418) and (hState = 552)) or
								((vState = 418) and (hState = 561)) or
								((vState = 418) and (hState = 562)) or
								((vState = 418) and (hState = 567)) or
								((vState = 418) and (hState = 588)) or
								((vState = 419) and (hState = 278)) or
								((vState = 419) and (hState = 279)) or
								((vState = 419) and (hState = 294)) or
								((vState = 419) and (hState = 298)) or
								((vState = 419) and (hState = 299)) or
								((vState = 419) and (hState = 310)) or
								((vState = 419) and (hState = 330)) or
								((vState = 419) and (hState = 331)) or
								((vState = 419) and (hState = 335)) or
								((vState = 419) and (hState = 345)) or
								((vState = 419) and (hState = 346)) or
								((vState = 419) and (hState = 347)) or
								((vState = 419) and (hState = 362)) or
								((vState = 419) and (hState = 382)) or
								((vState = 419) and (hState = 390)) or
								((vState = 419) and (hState = 396)) or
								((vState = 419) and (hState = 437)) or
								((vState = 419) and (hState = 438)) or
								((vState = 419) and (hState = 439)) or
								((vState = 419) and (hState = 440)) or
								((vState = 419) and (hState = 441)) or
								((vState = 419) and (hState = 442)) or
								((vState = 419) and (hState = 443)) or
								((vState = 419) and (hState = 444)) or
								((vState = 419) and (hState = 445)) or
								((vState = 419) and (hState = 469)) or
								((vState = 419) and (hState = 485)) or
								((vState = 419) and (hState = 501)) or
								((vState = 419) and (hState = 502)) or
								((vState = 419) and (hState = 511)) or
								((vState = 419) and (hState = 522)) or
								((vState = 419) and (hState = 529)) or
								((vState = 419) and (hState = 530)) or
								((vState = 419) and (hState = 531)) or
								((vState = 419) and (hState = 532)) or
								((vState = 419) and (hState = 533)) or
								((vState = 419) and (hState = 534)) or
								((vState = 419) and (hState = 535)) or
								((vState = 419) and (hState = 547)) or
								((vState = 419) and (hState = 548)) or
								((vState = 419) and (hState = 552)) or
								((vState = 419) and (hState = 560)) or
								((vState = 419) and (hState = 561)) or
								((vState = 419) and (hState = 567)) or
								((vState = 419) and (hState = 588)) or
								((vState = 420) and (hState = 294)) or
								((vState = 420) and (hState = 298)) or
								((vState = 420) and (hState = 299)) or
								((vState = 420) and (hState = 335)) or
								((vState = 420) and (hState = 345)) or
								((vState = 420) and (hState = 346)) or
								((vState = 420) and (hState = 361)) or
								((vState = 420) and (hState = 381)) or
								((vState = 420) and (hState = 382)) or
								((vState = 420) and (hState = 391)) or
								((vState = 420) and (hState = 396)) or
								((vState = 420) and (hState = 436)) or
								((vState = 420) and (hState = 437)) or
								((vState = 420) and (hState = 443)) or
								((vState = 420) and (hState = 444)) or
								((vState = 420) and (hState = 469)) or
								((vState = 420) and (hState = 485)) or
								((vState = 420) and (hState = 522)) or
								((vState = 420) and (hState = 529)) or
								((vState = 420) and (hState = 530)) or
								((vState = 420) and (hState = 531)) or
								((vState = 420) and (hState = 532)) or
								((vState = 420) and (hState = 533)) or
								((vState = 420) and (hState = 534)) or
								((vState = 420) and (hState = 535)) or
								((vState = 420) and (hState = 547)) or
								((vState = 420) and (hState = 548)) or
								((vState = 420) and (hState = 549)) or
								((vState = 420) and (hState = 560)) or
								((vState = 420) and (hState = 567)) or
								((vState = 420) and (hState = 588)) or
								((vState = 421) and (hState = 275)) or
								((vState = 421) and (hState = 298)) or
								((vState = 421) and (hState = 299)) or
								((vState = 421) and (hState = 321)) or
								((vState = 421) and (hState = 322)) or
								((vState = 421) and (hState = 335)) or
								((vState = 421) and (hState = 345)) or
								((vState = 421) and (hState = 346)) or
								((vState = 421) and (hState = 380)) or
								((vState = 421) and (hState = 381)) or
								((vState = 421) and (hState = 382)) or
								((vState = 421) and (hState = 392)) or
								((vState = 421) and (hState = 396)) or
								((vState = 421) and (hState = 419)) or
								((vState = 421) and (hState = 420)) or
								((vState = 421) and (hState = 437)) or
								((vState = 421) and (hState = 443)) or
								((vState = 421) and (hState = 469)) or
								((vState = 421) and (hState = 485)) or
								((vState = 421) and (hState = 503)) or
								((vState = 421) and (hState = 522)) or
								((vState = 421) and (hState = 529)) or
								((vState = 421) and (hState = 530)) or
								((vState = 421) and (hState = 535)) or
								((vState = 421) and (hState = 536)) or
								((vState = 421) and (hState = 538)) or
								((vState = 421) and (hState = 547)) or
								((vState = 421) and (hState = 548)) or
								((vState = 421) and (hState = 549)) or
								((vState = 421) and (hState = 560)) or
								((vState = 421) and (hState = 588)) or
								((vState = 422) and (hState = 297)) or
								((vState = 422) and (hState = 298)) or
								((vState = 422) and (hState = 299)) or
								((vState = 422) and (hState = 309)) or
								((vState = 422) and (hState = 319)) or
								((vState = 422) and (hState = 320)) or
								((vState = 422) and (hState = 321)) or
								((vState = 422) and (hState = 322)) or
								((vState = 422) and (hState = 323)) or
								((vState = 422) and (hState = 324)) or
								((vState = 422) and (hState = 335)) or
								((vState = 422) and (hState = 345)) or
								((vState = 422) and (hState = 346)) or
								((vState = 422) and (hState = 378)) or
								((vState = 422) and (hState = 379)) or
								((vState = 422) and (hState = 380)) or
								((vState = 422) and (hState = 381)) or
								((vState = 422) and (hState = 382)) or
								((vState = 422) and (hState = 392)) or
								((vState = 422) and (hState = 393)) or
								((vState = 422) and (hState = 396)) or
								((vState = 422) and (hState = 418)) or
								((vState = 422) and (hState = 419)) or
								((vState = 422) and (hState = 420)) or
								((vState = 422) and (hState = 421)) or
								((vState = 422) and (hState = 422)) or
								((vState = 422) and (hState = 423)) or
								((vState = 422) and (hState = 424)) or
								((vState = 422) and (hState = 437)) or
								((vState = 422) and (hState = 443)) or
								((vState = 422) and (hState = 459)) or
								((vState = 422) and (hState = 469)) or
								((vState = 422) and (hState = 485)) or
								((vState = 422) and (hState = 495)) or
								((vState = 422) and (hState = 496)) or
								((vState = 422) and (hState = 497)) or
								((vState = 422) and (hState = 503)) or
								((vState = 422) and (hState = 508)) or
								((vState = 422) and (hState = 529)) or
								((vState = 422) and (hState = 530)) or
								((vState = 422) and (hState = 535)) or
								((vState = 422) and (hState = 536)) or
								((vState = 422) and (hState = 537)) or
								((vState = 422) and (hState = 538)) or
								((vState = 422) and (hState = 547)) or
								((vState = 422) and (hState = 548)) or
								((vState = 422) and (hState = 560)) or
								((vState = 422) and (hState = 588)) or
								((vState = 422) and (hState = 593)) or
								((vState = 423) and (hState = 265)) or
								((vState = 423) and (hState = 273)) or
								((vState = 423) and (hState = 293)) or
								((vState = 423) and (hState = 297)) or
								((vState = 423) and (hState = 298)) or
								((vState = 423) and (hState = 299)) or
								((vState = 423) and (hState = 300)) or
								((vState = 423) and (hState = 309)) or
								((vState = 423) and (hState = 319)) or
								((vState = 423) and (hState = 320)) or
								((vState = 423) and (hState = 336)) or
								((vState = 423) and (hState = 345)) or
								((vState = 423) and (hState = 346)) or
								((vState = 423) and (hState = 378)) or
								((vState = 423) and (hState = 379)) or
								((vState = 423) and (hState = 380)) or
								((vState = 423) and (hState = 381)) or
								((vState = 423) and (hState = 382)) or
								((vState = 423) and (hState = 383)) or
								((vState = 423) and (hState = 394)) or
								((vState = 423) and (hState = 395)) or
								((vState = 423) and (hState = 396)) or
								((vState = 423) and (hState = 397)) or
								((vState = 423) and (hState = 398)) or
								((vState = 423) and (hState = 399)) or
								((vState = 423) and (hState = 400)) or
								((vState = 423) and (hState = 401)) or
								((vState = 423) and (hState = 402)) or
								((vState = 423) and (hState = 403)) or
								((vState = 423) and (hState = 404)) or
								((vState = 423) and (hState = 405)) or
								((vState = 423) and (hState = 406)) or
								((vState = 423) and (hState = 407)) or
								((vState = 423) and (hState = 408)) or
								((vState = 423) and (hState = 409)) or
								((vState = 423) and (hState = 410)) or
								((vState = 423) and (hState = 411)) or
								((vState = 423) and (hState = 412)) or
								((vState = 423) and (hState = 413)) or
								((vState = 423) and (hState = 414)) or
								((vState = 423) and (hState = 415)) or
								((vState = 423) and (hState = 416)) or
								((vState = 423) and (hState = 417)) or
								((vState = 423) and (hState = 418)) or
								((vState = 423) and (hState = 419)) or
								((vState = 423) and (hState = 420)) or
								((vState = 423) and (hState = 421)) or
								((vState = 423) and (hState = 422)) or
								((vState = 423) and (hState = 437)) or
								((vState = 423) and (hState = 469)) or
								((vState = 423) and (hState = 495)) or
								((vState = 423) and (hState = 496)) or
								((vState = 423) and (hState = 497)) or
								((vState = 423) and (hState = 505)) or
								((vState = 423) and (hState = 506)) or
								((vState = 423) and (hState = 529)) or
								((vState = 423) and (hState = 536)) or
								((vState = 423) and (hState = 537)) or
								((vState = 423) and (hState = 546)) or
								((vState = 423) and (hState = 547)) or
								((vState = 423) and (hState = 558)) or
								((vState = 423) and (hState = 559)) or
								((vState = 423) and (hState = 560)) or
								((vState = 423) and (hState = 568)) or
								((vState = 423) and (hState = 588)) or
								((vState = 423) and (hState = 593)) or
								((vState = 424) and (hState = 266)) or
								((vState = 424) and (hState = 272)) or
								((vState = 424) and (hState = 288)) or
								((vState = 424) and (hState = 293)) or
								((vState = 424) and (hState = 297)) or
								((vState = 424) and (hState = 298)) or
								((vState = 424) and (hState = 309)) or
								((vState = 424) and (hState = 320)) or
								((vState = 424) and (hState = 336)) or
								((vState = 424) and (hState = 345)) or
								((vState = 424) and (hState = 346)) or
								((vState = 424) and (hState = 377)) or
								((vState = 424) and (hState = 382)) or
								((vState = 424) and (hState = 383)) or
								((vState = 424) and (hState = 384)) or
								((vState = 424) and (hState = 409)) or
								((vState = 424) and (hState = 410)) or
								((vState = 424) and (hState = 411)) or
								((vState = 424) and (hState = 412)) or
								((vState = 424) and (hState = 413)) or
								((vState = 424) and (hState = 414)) or
								((vState = 424) and (hState = 415)) or
								((vState = 424) and (hState = 416)) or
								((vState = 424) and (hState = 417)) or
								((vState = 424) and (hState = 418)) or
								((vState = 424) and (hState = 419)) or
								((vState = 424) and (hState = 420)) or
								((vState = 424) and (hState = 421)) or
								((vState = 424) and (hState = 422)) or
								((vState = 424) and (hState = 437)) or
								((vState = 424) and (hState = 460)) or
								((vState = 424) and (hState = 486)) or
								((vState = 424) and (hState = 497)) or
								((vState = 424) and (hState = 505)) or
								((vState = 424) and (hState = 506)) or
								((vState = 424) and (hState = 523)) or
								((vState = 424) and (hState = 528)) or
								((vState = 424) and (hState = 529)) or
								((vState = 424) and (hState = 536)) or
								((vState = 424) and (hState = 545)) or
								((vState = 424) and (hState = 546)) or
								((vState = 424) and (hState = 547)) or
								((vState = 424) and (hState = 558)) or
								((vState = 424) and (hState = 559)) or
								((vState = 424) and (hState = 568)) or
								((vState = 424) and (hState = 588)) or
								((vState = 424) and (hState = 593)) or
								((vState = 425) and (hState = 287)) or
								((vState = 425) and (hState = 293)) or
								((vState = 425) and (hState = 297)) or
								((vState = 425) and (hState = 298)) or
								((vState = 425) and (hState = 302)) or
								((vState = 425) and (hState = 303)) or
								((vState = 425) and (hState = 304)) or
								((vState = 425) and (hState = 305)) or
								((vState = 425) and (hState = 345)) or
								((vState = 425) and (hState = 346)) or
								((vState = 425) and (hState = 356)) or
								((vState = 425) and (hState = 383)) or
								((vState = 425) and (hState = 384)) or
								((vState = 425) and (hState = 385)) or
								((vState = 425) and (hState = 415)) or
								((vState = 425) and (hState = 416)) or
								((vState = 425) and (hState = 417)) or
								((vState = 425) and (hState = 418)) or
								((vState = 425) and (hState = 419)) or
								((vState = 425) and (hState = 420)) or
								((vState = 425) and (hState = 421)) or
								((vState = 425) and (hState = 422)) or
								((vState = 425) and (hState = 423)) or
								((vState = 425) and (hState = 424)) or
								((vState = 425) and (hState = 425)) or
								((vState = 425) and (hState = 426)) or
								((vState = 425) and (hState = 427)) or
								((vState = 425) and (hState = 428)) or
								((vState = 425) and (hState = 429)) or
								((vState = 425) and (hState = 430)) or
								((vState = 425) and (hState = 431)) or
								((vState = 425) and (hState = 432)) or
								((vState = 425) and (hState = 433)) or
								((vState = 425) and (hState = 434)) or
								((vState = 425) and (hState = 435)) or
								((vState = 425) and (hState = 436)) or
								((vState = 425) and (hState = 437)) or
								((vState = 425) and (hState = 438)) or
								((vState = 425) and (hState = 439)) or
								((vState = 425) and (hState = 440)) or
								((vState = 425) and (hState = 487)) or
								((vState = 425) and (hState = 491)) or
								((vState = 425) and (hState = 503)) or
								((vState = 425) and (hState = 523)) or
								((vState = 425) and (hState = 527)) or
								((vState = 425) and (hState = 528)) or
								((vState = 425) and (hState = 529)) or
								((vState = 425) and (hState = 544)) or
								((vState = 425) and (hState = 545)) or
								((vState = 425) and (hState = 546)) or
								((vState = 425) and (hState = 547)) or
								((vState = 425) and (hState = 557)) or
								((vState = 425) and (hState = 558)) or
								((vState = 425) and (hState = 559)) or
								((vState = 425) and (hState = 568)) or
								((vState = 425) and (hState = 588)) or
								((vState = 426) and (hState = 267)) or
								((vState = 426) and (hState = 268)) or
								((vState = 426) and (hState = 269)) or
								((vState = 426) and (hState = 286)) or
								((vState = 426) and (hState = 293)) or
								((vState = 426) and (hState = 297)) or
								((vState = 426) and (hState = 298)) or
								((vState = 426) and (hState = 299)) or
								((vState = 426) and (hState = 300)) or
								((vState = 426) and (hState = 301)) or
								((vState = 426) and (hState = 302)) or
								((vState = 426) and (hState = 303)) or
								((vState = 426) and (hState = 304)) or
								((vState = 426) and (hState = 305)) or
								((vState = 426) and (hState = 306)) or
								((vState = 426) and (hState = 307)) or
								((vState = 426) and (hState = 308)) or
								((vState = 426) and (hState = 355)) or
								((vState = 426) and (hState = 373)) or
								((vState = 426) and (hState = 384)) or
								((vState = 426) and (hState = 385)) or
								((vState = 426) and (hState = 397)) or
								((vState = 426) and (hState = 415)) or
								((vState = 426) and (hState = 416)) or
								((vState = 426) and (hState = 417)) or
								((vState = 426) and (hState = 421)) or
								((vState = 426) and (hState = 422)) or
								((vState = 426) and (hState = 423)) or
								((vState = 426) and (hState = 424)) or
								((vState = 426) and (hState = 425)) or
								((vState = 426) and (hState = 426)) or
								((vState = 426) and (hState = 427)) or
								((vState = 426) and (hState = 428)) or
								((vState = 426) and (hState = 429)) or
								((vState = 426) and (hState = 430)) or
								((vState = 426) and (hState = 431)) or
								((vState = 426) and (hState = 432)) or
								((vState = 426) and (hState = 466)) or
								((vState = 426) and (hState = 487)) or
								((vState = 426) and (hState = 488)) or
								((vState = 426) and (hState = 489)) or
								((vState = 426) and (hState = 490)) or
								((vState = 426) and (hState = 502)) or
								((vState = 426) and (hState = 507)) or
								((vState = 426) and (hState = 523)) or
								((vState = 426) and (hState = 524)) or
								((vState = 426) and (hState = 525)) or
								((vState = 426) and (hState = 529)) or
								((vState = 426) and (hState = 537)) or
								((vState = 426) and (hState = 541)) or
								((vState = 426) and (hState = 545)) or
								((vState = 426) and (hState = 546)) or
								((vState = 426) and (hState = 547)) or
								((vState = 426) and (hState = 557)) or
								((vState = 426) and (hState = 558)) or
								((vState = 426) and (hState = 559)) or
								((vState = 426) and (hState = 568)) or
								((vState = 426) and (hState = 594)) or
								((vState = 426) and (hState = 599)) or
								((vState = 427) and (hState = 267)) or
								((vState = 427) and (hState = 268)) or
								((vState = 427) and (hState = 293)) or
								((vState = 427) and (hState = 297)) or
								((vState = 427) and (hState = 298)) or
								((vState = 427) and (hState = 299)) or
								((vState = 427) and (hState = 300)) or
								((vState = 427) and (hState = 301)) or
								((vState = 427) and (hState = 302)) or
								((vState = 427) and (hState = 303)) or
								((vState = 427) and (hState = 304)) or
								((vState = 427) and (hState = 305)) or
								((vState = 427) and (hState = 306)) or
								((vState = 427) and (hState = 307)) or
								((vState = 427) and (hState = 308)) or
								((vState = 427) and (hState = 355)) or
								((vState = 427) and (hState = 373)) or
								((vState = 427) and (hState = 384)) or
								((vState = 427) and (hState = 385)) or
								((vState = 427) and (hState = 397)) or
								((vState = 427) and (hState = 415)) or
								((vState = 427) and (hState = 416)) or
								((vState = 427) and (hState = 417)) or
								((vState = 427) and (hState = 421)) or
								((vState = 427) and (hState = 422)) or
								((vState = 427) and (hState = 423)) or
								((vState = 427) and (hState = 424)) or
								((vState = 427) and (hState = 425)) or
								((vState = 427) and (hState = 426)) or
								((vState = 427) and (hState = 427)) or
								((vState = 427) and (hState = 428)) or
								((vState = 427) and (hState = 429)) or
								((vState = 427) and (hState = 430)) or
								((vState = 427) and (hState = 431)) or
								((vState = 427) and (hState = 432)) or
								((vState = 427) and (hState = 466)) or
								((vState = 427) and (hState = 487)) or
								((vState = 427) and (hState = 488)) or
								((vState = 427) and (hState = 489)) or
								((vState = 427) and (hState = 490)) or
								((vState = 427) and (hState = 502)) or
								((vState = 427) and (hState = 507)) or
								((vState = 427) and (hState = 523)) or
								((vState = 427) and (hState = 524)) or
								((vState = 427) and (hState = 525)) or
								((vState = 427) and (hState = 529)) or
								((vState = 427) and (hState = 537)) or
								((vState = 427) and (hState = 538)) or
								((vState = 427) and (hState = 541)) or
								((vState = 427) and (hState = 545)) or
								((vState = 427) and (hState = 546)) or
								((vState = 427) and (hState = 547)) or
								((vState = 427) and (hState = 557)) or
								((vState = 427) and (hState = 558)) or
								((vState = 427) and (hState = 559)) or
								((vState = 427) and (hState = 568)) or
								((vState = 427) and (hState = 594)) or
								((vState = 427) and (hState = 599)) or
								((vState = 428) and (hState = 267)) or
								((vState = 428) and (hState = 268)) or
								((vState = 428) and (hState = 293)) or
								((vState = 428) and (hState = 294)) or
								((vState = 428) and (hState = 295)) or
								((vState = 428) and (hState = 296)) or
								((vState = 428) and (hState = 297)) or
								((vState = 428) and (hState = 298)) or
								((vState = 428) and (hState = 304)) or
								((vState = 428) and (hState = 305)) or
								((vState = 428) and (hState = 306)) or
								((vState = 428) and (hState = 307)) or
								((vState = 428) and (hState = 308)) or
								((vState = 428) and (hState = 352)) or
								((vState = 428) and (hState = 372)) or
								((vState = 428) and (hState = 384)) or
								((vState = 428) and (hState = 385)) or
								((vState = 428) and (hState = 386)) or
								((vState = 428) and (hState = 387)) or
								((vState = 428) and (hState = 397)) or
								((vState = 428) and (hState = 417)) or
								((vState = 428) and (hState = 428)) or
								((vState = 428) and (hState = 429)) or
								((vState = 428) and (hState = 430)) or
								((vState = 428) and (hState = 431)) or
								((vState = 428) and (hState = 432)) or
								((vState = 428) and (hState = 466)) or
								((vState = 428) and (hState = 487)) or
								((vState = 428) and (hState = 488)) or
								((vState = 428) and (hState = 489)) or
								((vState = 428) and (hState = 490)) or
								((vState = 428) and (hState = 499)) or
								((vState = 428) and (hState = 500)) or
								((vState = 428) and (hState = 501)) or
								((vState = 428) and (hState = 508)) or
								((vState = 428) and (hState = 523)) or
								((vState = 428) and (hState = 524)) or
								((vState = 428) and (hState = 529)) or
								((vState = 428) and (hState = 537)) or
								((vState = 428) and (hState = 538)) or
								((vState = 428) and (hState = 539)) or
								((vState = 428) and (hState = 540)) or
								((vState = 428) and (hState = 545)) or
								((vState = 428) and (hState = 546)) or
								((vState = 428) and (hState = 547)) or
								((vState = 428) and (hState = 594)) or
								((vState = 428) and (hState = 599)) or
								((vState = 429) and (hState = 291)) or
								((vState = 429) and (hState = 292)) or
								((vState = 429) and (hState = 293)) or
								((vState = 429) and (hState = 294)) or
								((vState = 429) and (hState = 295)) or
								((vState = 429) and (hState = 296)) or
								((vState = 429) and (hState = 297)) or
								((vState = 429) and (hState = 298)) or
								((vState = 429) and (hState = 304)) or
								((vState = 429) and (hState = 305)) or
								((vState = 429) and (hState = 306)) or
								((vState = 429) and (hState = 307)) or
								((vState = 429) and (hState = 308)) or
								((vState = 429) and (hState = 350)) or
								((vState = 429) and (hState = 371)) or
								((vState = 429) and (hState = 384)) or
								((vState = 429) and (hState = 388)) or
								((vState = 429) and (hState = 389)) or
								((vState = 429) and (hState = 397)) or
								((vState = 429) and (hState = 413)) or
								((vState = 429) and (hState = 417)) or
								((vState = 429) and (hState = 434)) or
								((vState = 429) and (hState = 435)) or
								((vState = 429) and (hState = 436)) or
								((vState = 429) and (hState = 437)) or
								((vState = 429) and (hState = 438)) or
								((vState = 429) and (hState = 439)) or
								((vState = 429) and (hState = 464)) or
								((vState = 429) and (hState = 465)) or
								((vState = 429) and (hState = 486)) or
								((vState = 429) and (hState = 490)) or
								((vState = 429) and (hState = 499)) or
								((vState = 429) and (hState = 500)) or
								((vState = 429) and (hState = 501)) or
								((vState = 429) and (hState = 523)) or
								((vState = 429) and (hState = 524)) or
								((vState = 429) and (hState = 529)) or
								((vState = 429) and (hState = 537)) or
								((vState = 429) and (hState = 538)) or
								((vState = 429) and (hState = 539)) or
								((vState = 429) and (hState = 540)) or
								((vState = 429) and (hState = 545)) or
								((vState = 429) and (hState = 546)) or
								((vState = 429) and (hState = 556)) or
								((vState = 429) and (hState = 569)) or
								((vState = 429) and (hState = 594)) or
								((vState = 429) and (hState = 599)) or
								((vState = 430) and (hState = 283)) or
								((vState = 430) and (hState = 284)) or
								((vState = 430) and (hState = 285)) or
								((vState = 430) and (hState = 286)) or
								((vState = 430) and (hState = 287)) or
								((vState = 430) and (hState = 288)) or
								((vState = 430) and (hState = 293)) or
								((vState = 430) and (hState = 294)) or
								((vState = 430) and (hState = 295)) or
								((vState = 430) and (hState = 296)) or
								((vState = 430) and (hState = 297)) or
								((vState = 430) and (hState = 298)) or
								((vState = 430) and (hState = 306)) or
								((vState = 430) and (hState = 384)) or
								((vState = 430) and (hState = 389)) or
								((vState = 430) and (hState = 390)) or
								((vState = 430) and (hState = 397)) or
								((vState = 430) and (hState = 412)) or
								((vState = 430) and (hState = 417)) or
								((vState = 430) and (hState = 434)) or
								((vState = 430) and (hState = 442)) or
								((vState = 430) and (hState = 443)) or
								((vState = 430) and (hState = 444)) or
								((vState = 430) and (hState = 445)) or
								((vState = 430) and (hState = 464)) or
								((vState = 430) and (hState = 465)) or
								((vState = 430) and (hState = 491)) or
								((vState = 430) and (hState = 497)) or
								((vState = 430) and (hState = 502)) or
								((vState = 430) and (hState = 521)) or
								((vState = 430) and (hState = 522)) or
								((vState = 430) and (hState = 523)) or
								((vState = 430) and (hState = 536)) or
								((vState = 430) and (hState = 540)) or
								((vState = 430) and (hState = 545)) or
								((vState = 430) and (hState = 546)) or
								((vState = 430) and (hState = 556)) or
								((vState = 430) and (hState = 557)) or
								((vState = 430) and (hState = 558)) or
								((vState = 430) and (hState = 569)) or
								((vState = 430) and (hState = 599)) or
								((vState = 431) and (hState = 262)) or
								((vState = 431) and (hState = 281)) or
								((vState = 431) and (hState = 282)) or
								((vState = 431) and (hState = 283)) or
								((vState = 431) and (hState = 293)) or
								((vState = 431) and (hState = 294)) or
								((vState = 431) and (hState = 295)) or
								((vState = 431) and (hState = 296)) or
								((vState = 431) and (hState = 297)) or
								((vState = 431) and (hState = 298)) or
								((vState = 431) and (hState = 306)) or
								((vState = 431) and (hState = 324)) or
								((vState = 431) and (hState = 346)) or
								((vState = 431) and (hState = 368)) or
								((vState = 431) and (hState = 389)) or
								((vState = 431) and (hState = 390)) or
								((vState = 431) and (hState = 391)) or
								((vState = 431) and (hState = 392)) or
								((vState = 431) and (hState = 397)) or
								((vState = 431) and (hState = 411)) or
								((vState = 431) and (hState = 434)) or
								((vState = 431) and (hState = 448)) or
								((vState = 431) and (hState = 449)) or
								((vState = 431) and (hState = 450)) or
								((vState = 431) and (hState = 451)) or
								((vState = 431) and (hState = 452)) or
								((vState = 431) and (hState = 453)) or
								((vState = 431) and (hState = 464)) or
								((vState = 431) and (hState = 465)) or
								((vState = 431) and (hState = 492)) or
								((vState = 431) and (hState = 496)) or
								((vState = 431) and (hState = 502)) or
								((vState = 431) and (hState = 503)) or
								((vState = 431) and (hState = 511)) or
								((vState = 431) and (hState = 519)) or
								((vState = 431) and (hState = 520)) or
								((vState = 431) and (hState = 521)) or
								((vState = 431) and (hState = 522)) or
								((vState = 431) and (hState = 528)) or
								((vState = 431) and (hState = 534)) or
								((vState = 431) and (hState = 535)) or
								((vState = 431) and (hState = 545)) or
								((vState = 431) and (hState = 546)) or
								((vState = 431) and (hState = 558)) or
								((vState = 431) and (hState = 569)) or
								((vState = 431) and (hState = 570)) or
								((vState = 431) and (hState = 595)) or
								((vState = 432) and (hState = 262)) or
								((vState = 432) and (hState = 281)) or
								((vState = 432) and (hState = 293)) or
								((vState = 432) and (hState = 294)) or
								((vState = 432) and (hState = 295)) or
								((vState = 432) and (hState = 296)) or
								((vState = 432) and (hState = 297)) or
								((vState = 432) and (hState = 298)) or
								((vState = 432) and (hState = 305)) or
								((vState = 432) and (hState = 306)) or
								((vState = 432) and (hState = 390)) or
								((vState = 432) and (hState = 391)) or
								((vState = 432) and (hState = 393)) or
								((vState = 432) and (hState = 397)) or
								((vState = 432) and (hState = 411)) or
								((vState = 432) and (hState = 434)) or
								((vState = 432) and (hState = 464)) or
								((vState = 432) and (hState = 465)) or
								((vState = 432) and (hState = 482)) or
								((vState = 432) and (hState = 492)) or
								((vState = 432) and (hState = 496)) or
								((vState = 432) and (hState = 502)) or
								((vState = 432) and (hState = 503)) or
								((vState = 432) and (hState = 511)) or
								((vState = 432) and (hState = 519)) or
								((vState = 432) and (hState = 520)) or
								((vState = 432) and (hState = 521)) or
								((vState = 432) and (hState = 528)) or
								((vState = 432) and (hState = 545)) or
								((vState = 432) and (hState = 546)) or
								((vState = 432) and (hState = 558)) or
								((vState = 432) and (hState = 570)) or
								((vState = 432) and (hState = 571)) or
								((vState = 432) and (hState = 595)) or
								((vState = 433) and (hState = 271)) or
								((vState = 433) and (hState = 280)) or
								((vState = 433) and (hState = 281)) or
								((vState = 433) and (hState = 293)) or
								((vState = 433) and (hState = 294)) or
								((vState = 433) and (hState = 295)) or
								((vState = 433) and (hState = 297)) or
								((vState = 433) and (hState = 298)) or
								((vState = 433) and (hState = 304)) or
								((vState = 433) and (hState = 305)) or
								((vState = 433) and (hState = 306)) or
								((vState = 433) and (hState = 325)) or
								((vState = 433) and (hState = 340)) or
								((vState = 433) and (hState = 385)) or
								((vState = 433) and (hState = 397)) or
								((vState = 433) and (hState = 416)) or
								((vState = 433) and (hState = 434)) or
								((vState = 433) and (hState = 466)) or
								((vState = 433) and (hState = 492)) or
								((vState = 433) and (hState = 493)) or
								((vState = 433) and (hState = 494)) or
								((vState = 433) and (hState = 495)) or
								((vState = 433) and (hState = 496)) or
								((vState = 433) and (hState = 504)) or
								((vState = 433) and (hState = 512)) or
								((vState = 433) and (hState = 518)) or
								((vState = 433) and (hState = 519)) or
								((vState = 433) and (hState = 520)) or
								((vState = 433) and (hState = 528)) or
								((vState = 433) and (hState = 532)) or
								((vState = 433) and (hState = 542)) or
								((vState = 433) and (hState = 543)) or
								((vState = 433) and (hState = 544)) or
								((vState = 433) and (hState = 545)) or
								((vState = 433) and (hState = 558)) or
								((vState = 433) and (hState = 571)) or
								((vState = 433) and (hState = 572)) or
								((vState = 433) and (hState = 585)) or
								((vState = 433) and (hState = 595)) or
								((vState = 434) and (hState = 271)) or
								((vState = 434) and (hState = 272)) or
								((vState = 434) and (hState = 273)) or
								((vState = 434) and (hState = 274)) or
								((vState = 434) and (hState = 281)) or
								((vState = 434) and (hState = 293)) or
								((vState = 434) and (hState = 294)) or
								((vState = 434) and (hState = 298)) or
								((vState = 434) and (hState = 304)) or
								((vState = 434) and (hState = 305)) or
								((vState = 434) and (hState = 306)) or
								((vState = 434) and (hState = 307)) or
								((vState = 434) and (hState = 308)) or
								((vState = 434) and (hState = 325)) or
								((vState = 434) and (hState = 340)) or
								((vState = 434) and (hState = 341)) or
								((vState = 434) and (hState = 342)) or
								((vState = 434) and (hState = 366)) or
								((vState = 434) and (hState = 385)) or
								((vState = 434) and (hState = 396)) or
								((vState = 434) and (hState = 397)) or
								((vState = 434) and (hState = 416)) or
								((vState = 434) and (hState = 434)) or
								((vState = 434) and (hState = 455)) or
								((vState = 434) and (hState = 466)) or
								((vState = 434) and (hState = 492)) or
								((vState = 434) and (hState = 493)) or
								((vState = 434) and (hState = 494)) or
								((vState = 434) and (hState = 495)) or
								((vState = 434) and (hState = 496)) or
								((vState = 434) and (hState = 497)) or
								((vState = 434) and (hState = 513)) or
								((vState = 434) and (hState = 517)) or
								((vState = 434) and (hState = 518)) or
								((vState = 434) and (hState = 519)) or
								((vState = 434) and (hState = 528)) or
								((vState = 434) and (hState = 529)) or
								((vState = 434) and (hState = 530)) or
								((vState = 434) and (hState = 531)) or
								((vState = 434) and (hState = 542)) or
								((vState = 434) and (hState = 543)) or
								((vState = 434) and (hState = 544)) or
								((vState = 434) and (hState = 545)) or
								((vState = 434) and (hState = 555)) or
								((vState = 434) and (hState = 556)) or
								((vState = 434) and (hState = 557)) or
								((vState = 434) and (hState = 571)) or
								((vState = 434) and (hState = 572)) or
								((vState = 434) and (hState = 573)) or
								((vState = 434) and (hState = 585)) or
								((vState = 434) and (hState = 595)) or
								((vState = 434) and (hState = 596)) or
								((vState = 434) and (hState = 597)) or
								((vState = 435) and (hState = 257)) or
								((vState = 435) and (hState = 269)) or
								((vState = 435) and (hState = 270)) or
								((vState = 435) and (hState = 271)) or
								((vState = 435) and (hState = 272)) or
								((vState = 435) and (hState = 293)) or
								((vState = 435) and (hState = 294)) or
								((vState = 435) and (hState = 298)) or
								((vState = 435) and (hState = 304)) or
								((vState = 435) and (hState = 305)) or
								((vState = 435) and (hState = 309)) or
								((vState = 435) and (hState = 326)) or
								((vState = 435) and (hState = 340)) or
								((vState = 435) and (hState = 341)) or
								((vState = 435) and (hState = 363)) or
								((vState = 435) and (hState = 385)) or
								((vState = 435) and (hState = 391)) or
								((vState = 435) and (hState = 397)) or
								((vState = 435) and (hState = 416)) or
								((vState = 435) and (hState = 489)) or
								((vState = 435) and (hState = 490)) or
								((vState = 435) and (hState = 491)) or
								((vState = 435) and (hState = 495)) or
								((vState = 435) and (hState = 496)) or
								((vState = 435) and (hState = 505)) or
								((vState = 435) and (hState = 506)) or
								((vState = 435) and (hState = 514)) or
								((vState = 435) and (hState = 515)) or
								((vState = 435) and (hState = 516)) or
								((vState = 435) and (hState = 517)) or
								((vState = 435) and (hState = 518)) or
								((vState = 435) and (hState = 528)) or
								((vState = 435) and (hState = 529)) or
								((vState = 435) and (hState = 542)) or
								((vState = 435) and (hState = 543)) or
								((vState = 435) and (hState = 544)) or
								((vState = 435) and (hState = 553)) or
								((vState = 435) and (hState = 554)) or
								((vState = 435) and (hState = 571)) or
								((vState = 435) and (hState = 572)) or
								((vState = 435) and (hState = 573)) or
								((vState = 435) and (hState = 574)) or
								((vState = 435) and (hState = 585)) or
								((vState = 435) and (hState = 597)) or
								((vState = 436) and (hState = 256)) or
								((vState = 436) and (hState = 265)) or
								((vState = 436) and (hState = 266)) or
								((vState = 436) and (hState = 272)) or
								((vState = 436) and (hState = 294)) or
								((vState = 436) and (hState = 298)) or
								((vState = 436) and (hState = 304)) or
								((vState = 436) and (hState = 305)) or
								((vState = 436) and (hState = 319)) or
								((vState = 436) and (hState = 326)) or
								((vState = 436) and (hState = 339)) or
								((vState = 436) and (hState = 340)) or
								((vState = 436) and (hState = 341)) or
								((vState = 436) and (hState = 362)) or
								((vState = 436) and (hState = 385)) or
								((vState = 436) and (hState = 392)) or
								((vState = 436) and (hState = 397)) or
								((vState = 436) and (hState = 398)) or
								((vState = 436) and (hState = 433)) or
								((vState = 436) and (hState = 469)) or
								((vState = 436) and (hState = 475)) or
								((vState = 436) and (hState = 476)) or
								((vState = 436) and (hState = 477)) or
								((vState = 436) and (hState = 484)) or
								((vState = 436) and (hState = 485)) or
								((vState = 436) and (hState = 486)) or
								((vState = 436) and (hState = 490)) or
								((vState = 436) and (hState = 491)) or
								((vState = 436) and (hState = 496)) or
								((vState = 436) and (hState = 505)) or
								((vState = 436) and (hState = 506)) or
								((vState = 436) and (hState = 507)) or
								((vState = 436) and (hState = 515)) or
								((vState = 436) and (hState = 516)) or
								((vState = 436) and (hState = 517)) or
								((vState = 436) and (hState = 528)) or
								((vState = 436) and (hState = 544)) or
								((vState = 436) and (hState = 552)) or
								((vState = 436) and (hState = 553)) or
								((vState = 436) and (hState = 571)) or
								((vState = 436) and (hState = 572)) or
								((vState = 436) and (hState = 585)) or
								((vState = 436) and (hState = 597)) or
								((vState = 437) and (hState = 255)) or
								((vState = 437) and (hState = 256)) or
								((vState = 437) and (hState = 273)) or
								((vState = 437) and (hState = 294)) or
								((vState = 437) and (hState = 298)) or
								((vState = 437) and (hState = 304)) or
								((vState = 437) and (hState = 305)) or
								((vState = 437) and (hState = 310)) or
								((vState = 437) and (hState = 319)) or
								((vState = 437) and (hState = 327)) or
								((vState = 437) and (hState = 361)) or
								((vState = 437) and (hState = 385)) or
								((vState = 437) and (hState = 386)) or
								((vState = 437) and (hState = 397)) or
								((vState = 437) and (hState = 398)) or
								((vState = 437) and (hState = 408)) or
								((vState = 437) and (hState = 433)) or
								((vState = 437) and (hState = 461)) or
								((vState = 437) and (hState = 469)) or
								((vState = 437) and (hState = 474)) or
								((vState = 437) and (hState = 475)) or
								((vState = 437) and (hState = 476)) or
								((vState = 437) and (hState = 477)) or
								((vState = 437) and (hState = 478)) or
								((vState = 437) and (hState = 490)) or
								((vState = 437) and (hState = 505)) or
								((vState = 437) and (hState = 506)) or
								((vState = 437) and (hState = 507)) or
								((vState = 437) and (hState = 513)) or
								((vState = 437) and (hState = 514)) or
								((vState = 437) and (hState = 515)) or
								((vState = 437) and (hState = 516)) or
								((vState = 437) and (hState = 517)) or
								((vState = 437) and (hState = 527)) or
								((vState = 437) and (hState = 528)) or
								((vState = 437) and (hState = 551)) or
								((vState = 437) and (hState = 552)) or
								((vState = 437) and (hState = 553)) or
								((vState = 437) and (hState = 571)) or
								((vState = 437) and (hState = 572)) or
								((vState = 437) and (hState = 585)) or
								((vState = 437) and (hState = 597)) or
								((vState = 438) and (hState = 255)) or
								((vState = 438) and (hState = 256)) or
								((vState = 438) and (hState = 294)) or
								((vState = 438) and (hState = 304)) or
								((vState = 438) and (hState = 305)) or
								((vState = 438) and (hState = 319)) or
								((vState = 438) and (hState = 385)) or
								((vState = 438) and (hState = 386)) or
								((vState = 438) and (hState = 387)) or
								((vState = 438) and (hState = 397)) or
								((vState = 438) and (hState = 433)) or
								((vState = 438) and (hState = 460)) or
								((vState = 438) and (hState = 461)) or
								((vState = 438) and (hState = 469)) or
								((vState = 438) and (hState = 474)) or
								((vState = 438) and (hState = 475)) or
								((vState = 438) and (hState = 490)) or
								((vState = 438) and (hState = 506)) or
								((vState = 438) and (hState = 507)) or
								((vState = 438) and (hState = 512)) or
								((vState = 438) and (hState = 513)) or
								((vState = 438) and (hState = 516)) or
								((vState = 438) and (hState = 517)) or
								((vState = 438) and (hState = 527)) or
								((vState = 438) and (hState = 528)) or
								((vState = 438) and (hState = 552)) or
								((vState = 438) and (hState = 572)) or
								((vState = 438) and (hState = 584)) or
								((vState = 438) and (hState = 597)) or
								((vState = 439) and (hState = 252)) or
								((vState = 439) and (hState = 253)) or
								((vState = 439) and (hState = 254)) or
								((vState = 439) and (hState = 255)) or
								((vState = 439) and (hState = 294)) or
								((vState = 439) and (hState = 303)) or
								((vState = 439) and (hState = 304)) or
								((vState = 439) and (hState = 305)) or
								((vState = 439) and (hState = 319)) or
								((vState = 439) and (hState = 320)) or
								((vState = 439) and (hState = 385)) or
								((vState = 439) and (hState = 386)) or
								((vState = 439) and (hState = 387)) or
								((vState = 439) and (hState = 397)) or
								((vState = 439) and (hState = 406)) or
								((vState = 439) and (hState = 433)) or
								((vState = 439) and (hState = 460)) or
								((vState = 439) and (hState = 461)) or
								((vState = 439) and (hState = 470)) or
								((vState = 439) and (hState = 471)) or
								((vState = 439) and (hState = 472)) or
								((vState = 439) and (hState = 506)) or
								((vState = 439) and (hState = 507)) or
								((vState = 439) and (hState = 508)) or
								((vState = 439) and (hState = 509)) or
								((vState = 439) and (hState = 510)) or
								((vState = 439) and (hState = 511)) or
								((vState = 439) and (hState = 512)) or
								((vState = 439) and (hState = 517)) or
								((vState = 439) and (hState = 528)) or
								((vState = 439) and (hState = 548)) or
								((vState = 439) and (hState = 552)) or
								((vState = 439) and (hState = 572)) or
								((vState = 439) and (hState = 584)) or
								((vState = 440) and (hState = 251)) or
								((vState = 440) and (hState = 252)) or
								((vState = 440) and (hState = 253)) or
								((vState = 440) and (hState = 254)) or
								((vState = 440) and (hState = 294)) or
								((vState = 440) and (hState = 303)) or
								((vState = 440) and (hState = 304)) or
								((vState = 440) and (hState = 319)) or
								((vState = 440) and (hState = 320)) or
								((vState = 440) and (hState = 321)) or
								((vState = 440) and (hState = 329)) or
								((vState = 440) and (hState = 384)) or
								((vState = 440) and (hState = 385)) or
								((vState = 440) and (hState = 386)) or
								((vState = 440) and (hState = 387)) or
								((vState = 440) and (hState = 395)) or
								((vState = 440) and (hState = 396)) or
								((vState = 440) and (hState = 405)) or
								((vState = 440) and (hState = 406)) or
								((vState = 440) and (hState = 460)) or
								((vState = 440) and (hState = 461)) or
								((vState = 440) and (hState = 462)) or
								((vState = 440) and (hState = 471)) or
								((vState = 440) and (hState = 506)) or
								((vState = 440) and (hState = 507)) or
								((vState = 440) and (hState = 508)) or
								((vState = 440) and (hState = 509)) or
								((vState = 440) and (hState = 510)) or
								((vState = 440) and (hState = 511)) or
								((vState = 440) and (hState = 512)) or
								((vState = 440) and (hState = 518)) or
								((vState = 440) and (hState = 522)) or
								((vState = 440) and (hState = 528)) or
								((vState = 440) and (hState = 547)) or
								((vState = 440) and (hState = 552)) or
								((vState = 440) and (hState = 572)) or
								((vState = 440) and (hState = 579)) or
								((vState = 440) and (hState = 583)) or
								((vState = 441) and (hState = 294)) or
								((vState = 441) and (hState = 295)) or
								((vState = 441) and (hState = 296)) or
								((vState = 441) and (hState = 297)) or
								((vState = 441) and (hState = 303)) or
								((vState = 441) and (hState = 304)) or
								((vState = 441) and (hState = 313)) or
								((vState = 441) and (hState = 319)) or
								((vState = 441) and (hState = 329)) or
								((vState = 441) and (hState = 330)) or
								((vState = 441) and (hState = 331)) or
								((vState = 441) and (hState = 383)) or
								((vState = 441) and (hState = 384)) or
								((vState = 441) and (hState = 385)) or
								((vState = 441) and (hState = 386)) or
								((vState = 441) and (hState = 387)) or
								((vState = 441) and (hState = 395)) or
								((vState = 441) and (hState = 396)) or
								((vState = 441) and (hState = 405)) or
								((vState = 441) and (hState = 406)) or
								((vState = 441) and (hState = 432)) or
								((vState = 441) and (hState = 459)) or
								((vState = 441) and (hState = 464)) or
								((vState = 441) and (hState = 471)) or
								((vState = 441) and (hState = 506)) or
								((vState = 441) and (hState = 507)) or
								((vState = 441) and (hState = 508)) or
								((vState = 441) and (hState = 509)) or
								((vState = 441) and (hState = 510)) or
								((vState = 441) and (hState = 511)) or
								((vState = 441) and (hState = 518)) or
								((vState = 441) and (hState = 519)) or
								((vState = 441) and (hState = 520)) or
								((vState = 441) and (hState = 544)) or
								((vState = 441) and (hState = 545)) or
								((vState = 441) and (hState = 551)) or
								((vState = 441) and (hState = 572)) or
								((vState = 441) and (hState = 581)) or
								((vState = 441) and (hState = 582)) or
								((vState = 441) and (hState = 583)) or
								((vState = 441) and (hState = 597)) or
								((vState = 442) and (hState = 276)) or
								((vState = 442) and (hState = 294)) or
								((vState = 442) and (hState = 295)) or
								((vState = 442) and (hState = 296)) or
								((vState = 442) and (hState = 297)) or
								((vState = 442) and (hState = 298)) or
								((vState = 442) and (hState = 299)) or
								((vState = 442) and (hState = 300)) or
								((vState = 442) and (hState = 301)) or
								((vState = 442) and (hState = 302)) or
								((vState = 442) and (hState = 303)) or
								((vState = 442) and (hState = 304)) or
								((vState = 442) and (hState = 314)) or
								((vState = 442) and (hState = 319)) or
								((vState = 442) and (hState = 329)) or
								((vState = 442) and (hState = 330)) or
								((vState = 442) and (hState = 331)) or
								((vState = 442) and (hState = 383)) or
								((vState = 442) and (hState = 384)) or
								((vState = 442) and (hState = 385)) or
								((vState = 442) and (hState = 386)) or
								((vState = 442) and (hState = 387)) or
								((vState = 442) and (hState = 388)) or
								((vState = 442) and (hState = 395)) or
								((vState = 442) and (hState = 396)) or
								((vState = 442) and (hState = 404)) or
								((vState = 442) and (hState = 408)) or
								((vState = 442) and (hState = 432)) or
								((vState = 442) and (hState = 459)) or
								((vState = 442) and (hState = 465)) or
								((vState = 442) and (hState = 487)) or
								((vState = 442) and (hState = 506)) or
								((vState = 442) and (hState = 507)) or
								((vState = 442) and (hState = 508)) or
								((vState = 442) and (hState = 509)) or
								((vState = 442) and (hState = 510)) or
								((vState = 442) and (hState = 511)) or
								((vState = 442) and (hState = 518)) or
								((vState = 442) and (hState = 519)) or
								((vState = 442) and (hState = 520)) or
								((vState = 442) and (hState = 527)) or
								((vState = 442) and (hState = 542)) or
								((vState = 442) and (hState = 543)) or
								((vState = 442) and (hState = 544)) or
								((vState = 442) and (hState = 551)) or
								((vState = 442) and (hState = 572)) or
								((vState = 442) and (hState = 582)) or
								((vState = 442) and (hState = 583)) or
								((vState = 442) and (hState = 597)) or
								((vState = 443) and (hState = 294)) or
								((vState = 443) and (hState = 295)) or
								((vState = 443) and (hState = 296)) or
								((vState = 443) and (hState = 297)) or
								((vState = 443) and (hState = 303)) or
								((vState = 443) and (hState = 304)) or
								((vState = 443) and (hState = 319)) or
								((vState = 443) and (hState = 331)) or
								((vState = 443) and (hState = 385)) or
								((vState = 443) and (hState = 386)) or
								((vState = 443) and (hState = 387)) or
								((vState = 443) and (hState = 388)) or
								((vState = 443) and (hState = 395)) or
								((vState = 443) and (hState = 396)) or
								((vState = 443) and (hState = 432)) or
								((vState = 443) and (hState = 487)) or
								((vState = 443) and (hState = 506)) or
								((vState = 443) and (hState = 507)) or
								((vState = 443) and (hState = 508)) or
								((vState = 443) and (hState = 511)) or
								((vState = 443) and (hState = 520)) or
								((vState = 443) and (hState = 527)) or
								((vState = 443) and (hState = 542)) or
								((vState = 443) and (hState = 543)) or
								((vState = 443) and (hState = 572)) or
								((vState = 443) and (hState = 582)) or
								((vState = 443) and (hState = 583)) or
								((vState = 443) and (hState = 597)) or
								((vState = 444) and (hState = 294)) or
								((vState = 444) and (hState = 295)) or
								((vState = 444) and (hState = 296)) or
								((vState = 444) and (hState = 297)) or
								((vState = 444) and (hState = 303)) or
								((vState = 444) and (hState = 304)) or
								((vState = 444) and (hState = 305)) or
								((vState = 444) and (hState = 319)) or
								((vState = 444) and (hState = 324)) or
								((vState = 444) and (hState = 331)) or
								((vState = 444) and (hState = 385)) or
								((vState = 444) and (hState = 386)) or
								((vState = 444) and (hState = 387)) or
								((vState = 444) and (hState = 388)) or
								((vState = 444) and (hState = 432)) or
								((vState = 444) and (hState = 501)) or
								((vState = 444) and (hState = 506)) or
								((vState = 444) and (hState = 507)) or
								((vState = 444) and (hState = 512)) or
								((vState = 444) and (hState = 527)) or
								((vState = 444) and (hState = 542)) or
								((vState = 444) and (hState = 597)) or
								((vState = 445) and (hState = 277)) or
								((vState = 445) and (hState = 294)) or
								((vState = 445) and (hState = 295)) or
								((vState = 445) and (hState = 296)) or
								((vState = 445) and (hState = 297)) or
								((vState = 445) and (hState = 303)) or
								((vState = 445) and (hState = 304)) or
								((vState = 445) and (hState = 308)) or
								((vState = 445) and (hState = 309)) or
								((vState = 445) and (hState = 315)) or
								((vState = 445) and (hState = 319)) or
								((vState = 445) and (hState = 324)) or
								((vState = 445) and (hState = 325)) or
								((vState = 445) and (hState = 331)) or
								((vState = 445) and (hState = 341)) or
								((vState = 445) and (hState = 385)) or
								((vState = 445) and (hState = 386)) or
								((vState = 445) and (hState = 387)) or
								((vState = 445) and (hState = 388)) or
								((vState = 445) and (hState = 402)) or
								((vState = 445) and (hState = 411)) or
								((vState = 445) and (hState = 432)) or
								((vState = 445) and (hState = 474)) or
								((vState = 445) and (hState = 486)) or
								((vState = 445) and (hState = 502)) or
								((vState = 445) and (hState = 503)) or
								((vState = 445) and (hState = 504)) or
								((vState = 445) and (hState = 505)) or
								((vState = 445) and (hState = 506)) or
								((vState = 445) and (hState = 507)) or
								((vState = 445) and (hState = 513)) or
								((vState = 445) and (hState = 514)) or
								((vState = 445) and (hState = 522)) or
								((vState = 445) and (hState = 527)) or
								((vState = 445) and (hState = 542)) or
								((vState = 445) and (hState = 584)) or
								((vState = 445) and (hState = 597)) or
								((vState = 446) and (hState = 278)) or
								((vState = 446) and (hState = 296)) or
								((vState = 446) and (hState = 297)) or
								((vState = 446) and (hState = 302)) or
								((vState = 446) and (hState = 303)) or
								((vState = 446) and (hState = 312)) or
								((vState = 446) and (hState = 313)) or
								((vState = 446) and (hState = 314)) or
								((vState = 446) and (hState = 315)) or
								((vState = 446) and (hState = 316)) or
								((vState = 446) and (hState = 317)) or
								((vState = 446) and (hState = 318)) or
								((vState = 446) and (hState = 319)) or
								((vState = 446) and (hState = 323)) or
								((vState = 446) and (hState = 324)) or
								((vState = 446) and (hState = 325)) or
								((vState = 446) and (hState = 341)) or
								((vState = 446) and (hState = 385)) or
								((vState = 446) and (hState = 400)) or
								((vState = 446) and (hState = 401)) or
								((vState = 446) and (hState = 413)) or
								((vState = 446) and (hState = 432)) or
								((vState = 446) and (hState = 433)) or
								((vState = 446) and (hState = 434)) or
								((vState = 446) and (hState = 435)) or
								((vState = 446) and (hState = 436)) or
								((vState = 446) and (hState = 437)) or
								((vState = 446) and (hState = 469)) or
								((vState = 446) and (hState = 475)) or
								((vState = 446) and (hState = 486)) or
								((vState = 446) and (hState = 502)) or
								((vState = 446) and (hState = 503)) or
								((vState = 446) and (hState = 504)) or
								((vState = 446) and (hState = 505)) or
								((vState = 446) and (hState = 506)) or
								((vState = 446) and (hState = 507)) or
								((vState = 446) and (hState = 536)) or
								((vState = 446) and (hState = 537)) or
								((vState = 446) and (hState = 542)) or
								((vState = 446) and (hState = 585)) or
								((vState = 446) and (hState = 597)) or
								((vState = 447) and (hState = 278)) or
								((vState = 447) and (hState = 296)) or
								((vState = 447) and (hState = 297)) or
								((vState = 447) and (hState = 302)) or
								((vState = 447) and (hState = 303)) or
								((vState = 447) and (hState = 315)) or
								((vState = 447) and (hState = 316)) or
								((vState = 447) and (hState = 317)) or
								((vState = 447) and (hState = 318)) or
								((vState = 447) and (hState = 319)) or
								((vState = 447) and (hState = 320)) or
								((vState = 447) and (hState = 321)) or
								((vState = 447) and (hState = 326)) or
								((vState = 447) and (hState = 379)) or
								((vState = 447) and (hState = 385)) or
								((vState = 447) and (hState = 389)) or
								((vState = 447) and (hState = 400)) or
								((vState = 447) and (hState = 401)) or
								((vState = 447) and (hState = 439)) or
								((vState = 447) and (hState = 440)) or
								((vState = 447) and (hState = 441)) or
								((vState = 447) and (hState = 442)) or
								((vState = 447) and (hState = 443)) or
								((vState = 447) and (hState = 470)) or
								((vState = 447) and (hState = 485)) or
								((vState = 447) and (hState = 501)) or
								((vState = 447) and (hState = 502)) or
								((vState = 447) and (hState = 503)) or
								((vState = 447) and (hState = 504)) or
								((vState = 447) and (hState = 505)) or
								((vState = 447) and (hState = 506)) or
								((vState = 447) and (hState = 507)) or
								((vState = 447) and (hState = 523)) or
								((vState = 447) and (hState = 524)) or
								((vState = 447) and (hState = 525)) or
								((vState = 447) and (hState = 535)) or
								((vState = 447) and (hState = 542)) or
								((vState = 447) and (hState = 579)) or
								((vState = 448) and (hState = 296)) or
								((vState = 448) and (hState = 297)) or
								((vState = 448) and (hState = 302)) or
								((vState = 448) and (hState = 303)) or
								((vState = 448) and (hState = 318)) or
								((vState = 448) and (hState = 319)) or
								((vState = 448) and (hState = 320)) or
								((vState = 448) and (hState = 321)) or
								((vState = 448) and (hState = 326)) or
								((vState = 448) and (hState = 385)) or
								((vState = 448) and (hState = 389)) or
								((vState = 448) and (hState = 400)) or
								((vState = 448) and (hState = 401)) or
								((vState = 448) and (hState = 439)) or
								((vState = 448) and (hState = 440)) or
								((vState = 448) and (hState = 441)) or
								((vState = 448) and (hState = 442)) or
								((vState = 448) and (hState = 443)) or
								((vState = 448) and (hState = 485)) or
								((vState = 448) and (hState = 501)) or
								((vState = 448) and (hState = 502)) or
								((vState = 448) and (hState = 503)) or
								((vState = 448) and (hState = 504)) or
								((vState = 448) and (hState = 505)) or
								((vState = 448) and (hState = 506)) or
								((vState = 448) and (hState = 507)) or
								((vState = 448) and (hState = 523)) or
								((vState = 448) and (hState = 524)) or
								((vState = 448) and (hState = 525)) or
								((vState = 448) and (hState = 535)) or
								((vState = 448) and (hState = 542)) or
								((vState = 448) and (hState = 579)) or
								((vState = 449) and (hState = 296)) or
								((vState = 449) and (hState = 297)) or
								((vState = 449) and (hState = 302)) or
								((vState = 449) and (hState = 303)) or
								((vState = 449) and (hState = 319)) or
								((vState = 449) and (hState = 326)) or
								((vState = 449) and (hState = 327)) or
								((vState = 449) and (hState = 340)) or
								((vState = 449) and (hState = 361)) or
								((vState = 449) and (hState = 385)) or
								((vState = 449) and (hState = 389)) or
								((vState = 449) and (hState = 392)) or
								((vState = 449) and (hState = 429)) or
								((vState = 449) and (hState = 430)) or
								((vState = 449) and (hState = 439)) or
								((vState = 449) and (hState = 440)) or
								((vState = 449) and (hState = 441)) or
								((vState = 449) and (hState = 442)) or
								((vState = 449) and (hState = 443)) or
								((vState = 449) and (hState = 444)) or
								((vState = 449) and (hState = 445)) or
								((vState = 449) and (hState = 446)) or
								((vState = 449) and (hState = 447)) or
								((vState = 449) and (hState = 448)) or
								((vState = 449) and (hState = 449)) or
								((vState = 449) and (hState = 455)) or
								((vState = 449) and (hState = 476)) or
								((vState = 449) and (hState = 501)) or
								((vState = 449) and (hState = 502)) or
								((vState = 449) and (hState = 505)) or
								((vState = 449) and (hState = 506)) or
								((vState = 449) and (hState = 507)) or
								((vState = 449) and (hState = 508)) or
								((vState = 449) and (hState = 525)) or
								((vState = 449) and (hState = 532)) or
								((vState = 449) and (hState = 533)) or
								((vState = 449) and (hState = 534)) or
								((vState = 449) and (hState = 535)) or
								((vState = 449) and (hState = 542)) or
								((vState = 449) and (hState = 548)) or
								((vState = 449) and (hState = 595)) or
								((vState = 450) and (hState = 281)) or
								((vState = 450) and (hState = 296)) or
								((vState = 450) and (hState = 297)) or
								((vState = 450) and (hState = 302)) or
								((vState = 450) and (hState = 303)) or
								((vState = 450) and (hState = 319)) or
								((vState = 450) and (hState = 324)) or
								((vState = 450) and (hState = 325)) or
								((vState = 450) and (hState = 326)) or
								((vState = 450) and (hState = 327)) or
								((vState = 450) and (hState = 340)) or
								((vState = 450) and (hState = 361)) or
								((vState = 450) and (hState = 378)) or
								((vState = 450) and (hState = 385)) or
								((vState = 450) and (hState = 389)) or
								((vState = 450) and (hState = 402)) or
								((vState = 450) and (hState = 421)) or
								((vState = 450) and (hState = 422)) or
								((vState = 450) and (hState = 423)) or
								((vState = 450) and (hState = 424)) or
								((vState = 450) and (hState = 425)) or
								((vState = 450) and (hState = 426)) or
								((vState = 450) and (hState = 427)) or
								((vState = 450) and (hState = 428)) or
								((vState = 450) and (hState = 429)) or
								((vState = 450) and (hState = 430)) or
								((vState = 450) and (hState = 431)) or
								((vState = 450) and (hState = 432)) or
								((vState = 450) and (hState = 433)) or
								((vState = 450) and (hState = 434)) or
								((vState = 450) and (hState = 435)) or
								((vState = 450) and (hState = 436)) or
								((vState = 450) and (hState = 437)) or
								((vState = 450) and (hState = 438)) or
								((vState = 450) and (hState = 439)) or
								((vState = 450) and (hState = 440)) or
								((vState = 450) and (hState = 441)) or
								((vState = 450) and (hState = 442)) or
								((vState = 450) and (hState = 443)) or
								((vState = 450) and (hState = 444)) or
								((vState = 450) and (hState = 445)) or
								((vState = 450) and (hState = 446)) or
								((vState = 450) and (hState = 447)) or
								((vState = 450) and (hState = 448)) or
								((vState = 450) and (hState = 449)) or
								((vState = 450) and (hState = 450)) or
								((vState = 450) and (hState = 451)) or
								((vState = 450) and (hState = 452)) or
								((vState = 450) and (hState = 453)) or
								((vState = 450) and (hState = 454)) or
								((vState = 450) and (hState = 455)) or
								((vState = 450) and (hState = 474)) or
								((vState = 450) and (hState = 475)) or
								((vState = 450) and (hState = 476)) or
								((vState = 450) and (hState = 477)) or
								((vState = 450) and (hState = 501)) or
								((vState = 450) and (hState = 502)) or
								((vState = 450) and (hState = 506)) or
								((vState = 450) and (hState = 507)) or
								((vState = 450) and (hState = 508)) or
								((vState = 450) and (hState = 525)) or
								((vState = 450) and (hState = 529)) or
								((vState = 450) and (hState = 530)) or
								((vState = 450) and (hState = 531)) or
								((vState = 450) and (hState = 532)) or
								((vState = 450) and (hState = 533)) or
								((vState = 450) and (hState = 534)) or
								((vState = 450) and (hState = 535)) or
								((vState = 450) and (hState = 536)) or
								((vState = 450) and (hState = 537)) or
								((vState = 450) and (hState = 538)) or
								((vState = 450) and (hState = 539)) or
								((vState = 450) and (hState = 540)) or
								((vState = 450) and (hState = 541)) or
								((vState = 450) and (hState = 542)) or
								((vState = 450) and (hState = 543)) or
								((vState = 450) and (hState = 544)) or
								((vState = 450) and (hState = 545)) or
								((vState = 450) and (hState = 546)) or
								((vState = 450) and (hState = 547)) or
								((vState = 450) and (hState = 548)) or
								((vState = 450) and (hState = 549)) or
								((vState = 450) and (hState = 550)) or
								((vState = 450) and (hState = 551)) or
								((vState = 450) and (hState = 552)) or
								((vState = 450) and (hState = 553)) or
								((vState = 450) and (hState = 578)) or
								((vState = 450) and (hState = 589)) or
								((vState = 450) and (hState = 595)) or
								((vState = 451) and (hState = 296)) or
								((vState = 451) and (hState = 297)) or
								((vState = 451) and (hState = 319)) or
								((vState = 451) and (hState = 328)) or
								((vState = 451) and (hState = 329)) or
								((vState = 451) and (hState = 330)) or
								((vState = 451) and (hState = 335)) or
								((vState = 451) and (hState = 361)) or
								((vState = 451) and (hState = 385)) or
								((vState = 451) and (hState = 390)) or
								((vState = 451) and (hState = 391)) or
								((vState = 451) and (hState = 426)) or
								((vState = 451) and (hState = 427)) or
								((vState = 451) and (hState = 428)) or
								((vState = 451) and (hState = 429)) or
								((vState = 451) and (hState = 454)) or
								((vState = 451) and (hState = 455)) or
								((vState = 451) and (hState = 456)) or
								((vState = 451) and (hState = 457)) or
								((vState = 451) and (hState = 458)) or
								((vState = 451) and (hState = 459)) or
								((vState = 451) and (hState = 460)) or
								((vState = 451) and (hState = 461)) or
								((vState = 451) and (hState = 475)) or
								((vState = 451) and (hState = 476)) or
								((vState = 451) and (hState = 477)) or
								((vState = 451) and (hState = 501)) or
								((vState = 451) and (hState = 507)) or
								((vState = 451) and (hState = 508)) or
								((vState = 451) and (hState = 525)) or
								((vState = 451) and (hState = 529)) or
								((vState = 451) and (hState = 539)) or
								((vState = 451) and (hState = 540)) or
								((vState = 451) and (hState = 545)) or
								((vState = 451) and (hState = 546)) or
								((vState = 451) and (hState = 547)) or
								((vState = 451) and (hState = 548)) or
								((vState = 451) and (hState = 549)) or
								((vState = 451) and (hState = 550)) or
								((vState = 451) and (hState = 551)) or
								((vState = 451) and (hState = 552)) or
								((vState = 451) and (hState = 553)) or
								((vState = 451) and (hState = 578)) or
								((vState = 451) and (hState = 590)) or
								((vState = 451) and (hState = 594)) or
								((vState = 451) and (hState = 595)) or
								((vState = 452) and (hState = 282)) or
								((vState = 452) and (hState = 296)) or
								((vState = 452) and (hState = 297)) or
								((vState = 452) and (hState = 301)) or
								((vState = 452) and (hState = 319)) or
								((vState = 452) and (hState = 330)) or
								((vState = 452) and (hState = 331)) or
								((vState = 452) and (hState = 332)) or
								((vState = 452) and (hState = 333)) or
								((vState = 452) and (hState = 334)) or
								((vState = 452) and (hState = 335)) or
								((vState = 452) and (hState = 361)) or
								((vState = 452) and (hState = 377)) or
								((vState = 452) and (hState = 385)) or
								((vState = 452) and (hState = 390)) or
								((vState = 452) and (hState = 391)) or
								((vState = 452) and (hState = 397)) or
								((vState = 452) and (hState = 429)) or
								((vState = 452) and (hState = 454)) or
								((vState = 452) and (hState = 462)) or
								((vState = 452) and (hState = 463)) or
								((vState = 452) and (hState = 464)) or
								((vState = 452) and (hState = 465)) or
								((vState = 452) and (hState = 466)) or
								((vState = 452) and (hState = 467)) or
								((vState = 452) and (hState = 476)) or
								((vState = 452) and (hState = 477)) or
								((vState = 452) and (hState = 478)) or
								((vState = 452) and (hState = 507)) or
								((vState = 452) and (hState = 508)) or
								((vState = 452) and (hState = 524)) or
								((vState = 452) and (hState = 525)) or
								((vState = 452) and (hState = 526)) or
								((vState = 452) and (hState = 527)) or
								((vState = 452) and (hState = 528)) or
								((vState = 452) and (hState = 539)) or
								((vState = 452) and (hState = 540)) or
								((vState = 452) and (hState = 545)) or
								((vState = 452) and (hState = 546)) or
								((vState = 452) and (hState = 547)) or
								((vState = 452) and (hState = 548)) or
								((vState = 452) and (hState = 577)) or
								((vState = 452) and (hState = 592)) or
								((vState = 452) and (hState = 593)) or
								((vState = 452) and (hState = 594)) or
								((vState = 452) and (hState = 595)) or
								((vState = 453) and (hState = 296)) or
								((vState = 453) and (hState = 297)) or
								((vState = 453) and (hState = 301)) or
								((vState = 453) and (hState = 319)) or
								((vState = 453) and (hState = 331)) or
								((vState = 453) and (hState = 361)) or
								((vState = 453) and (hState = 376)) or
								((vState = 453) and (hState = 385)) or
								((vState = 453) and (hState = 390)) or
								((vState = 453) and (hState = 429)) or
								((vState = 453) and (hState = 466)) or
								((vState = 453) and (hState = 467)) or
								((vState = 453) and (hState = 468)) or
								((vState = 453) and (hState = 477)) or
								((vState = 453) and (hState = 478)) or
								((vState = 453) and (hState = 479)) or
								((vState = 453) and (hState = 482)) or
								((vState = 453) and (hState = 508)) or
								((vState = 453) and (hState = 524)) or
								((vState = 453) and (hState = 525)) or
								((vState = 453) and (hState = 526)) or
								((vState = 453) and (hState = 527)) or
								((vState = 453) and (hState = 528)) or
								((vState = 453) and (hState = 539)) or
								((vState = 453) and (hState = 540)) or
								((vState = 453) and (hState = 546)) or
								((vState = 453) and (hState = 577)) or
								((vState = 453) and (hState = 592)) or
								((vState = 453) and (hState = 593)) or
								((vState = 453) and (hState = 594)) or
								((vState = 454) and (hState = 301)) or
								((vState = 454) and (hState = 319)) or
								((vState = 454) and (hState = 331)) or
								((vState = 454) and (hState = 337)) or
								((vState = 454) and (hState = 338)) or
								((vState = 454) and (hState = 361)) or
								((vState = 454) and (hState = 395)) or
								((vState = 454) and (hState = 396)) or
								((vState = 454) and (hState = 429)) or
								((vState = 454) and (hState = 453)) or
								((vState = 454) and (hState = 466)) or
								((vState = 454) and (hState = 478)) or
								((vState = 454) and (hState = 479)) or
								((vState = 454) and (hState = 480)) or
								((vState = 454) and (hState = 481)) or
								((vState = 454) and (hState = 509)) or
								((vState = 454) and (hState = 524)) or
								((vState = 454) and (hState = 537)) or
								((vState = 454) and (hState = 538)) or
								((vState = 454) and (hState = 546)) or
								((vState = 454) and (hState = 594)) or
								((vState = 455) and (hState = 301)) or
								((vState = 455) and (hState = 319)) or
								((vState = 455) and (hState = 338)) or
								((vState = 455) and (hState = 339)) or
								((vState = 455) and (hState = 361)) or
								((vState = 455) and (hState = 395)) or
								((vState = 455) and (hState = 396)) or
								((vState = 455) and (hState = 429)) or
								((vState = 455) and (hState = 466)) or
								((vState = 455) and (hState = 471)) or
								((vState = 455) and (hState = 472)) or
								((vState = 455) and (hState = 478)) or
								((vState = 455) and (hState = 479)) or
								((vState = 455) and (hState = 480)) or
								((vState = 455) and (hState = 481)) or
								((vState = 455) and (hState = 523)) or
								((vState = 455) and (hState = 524)) or
								((vState = 455) and (hState = 529)) or
								((vState = 455) and (hState = 534)) or
								((vState = 455) and (hState = 535)) or
								((vState = 455) and (hState = 536)) or
								((vState = 455) and (hState = 590)) or
								((vState = 455) and (hState = 594)) or
								((vState = 456) and (hState = 319)) or
								((vState = 456) and (hState = 338)) or
								((vState = 456) and (hState = 374)) or
								((vState = 456) and (hState = 389)) or
								((vState = 456) and (hState = 395)) or
								((vState = 456) and (hState = 396)) or
								((vState = 456) and (hState = 421)) or
								((vState = 456) and (hState = 429)) or
								((vState = 456) and (hState = 465)) or
								((vState = 456) and (hState = 466)) or
								((vState = 456) and (hState = 471)) or
								((vState = 456) and (hState = 472)) or
								((vState = 456) and (hState = 473)) or
								((vState = 456) and (hState = 474)) or
								((vState = 456) and (hState = 475)) or
								((vState = 456) and (hState = 476)) or
								((vState = 456) and (hState = 477)) or
								((vState = 456) and (hState = 478)) or
								((vState = 456) and (hState = 479)) or
								((vState = 456) and (hState = 480)) or
								((vState = 456) and (hState = 481)) or
								((vState = 456) and (hState = 521)) or
								((vState = 456) and (hState = 522)) or
								((vState = 456) and (hState = 523)) or
								((vState = 456) and (hState = 524)) or
								((vState = 456) and (hState = 529)) or
								((vState = 456) and (hState = 530)) or
								((vState = 456) and (hState = 531)) or
								((vState = 456) and (hState = 532)) or
								((vState = 456) and (hState = 533)) or
								((vState = 456) and (hState = 534)) or
								((vState = 456) and (hState = 535)) or
								((vState = 456) and (hState = 589)) or
								((vState = 456) and (hState = 594)) or
								((vState = 456) and (hState = 595)) or
								((vState = 457) and (hState = 319)) or
								((vState = 457) and (hState = 338)) or
								((vState = 457) and (hState = 346)) or
								((vState = 457) and (hState = 362)) or
								((vState = 457) and (hState = 373)) or
								((vState = 457) and (hState = 384)) or
								((vState = 457) and (hState = 394)) or
								((vState = 457) and (hState = 397)) or
								((vState = 457) and (hState = 463)) or
								((vState = 457) and (hState = 464)) or
								((vState = 457) and (hState = 465)) or
								((vState = 457) and (hState = 466)) or
								((vState = 457) and (hState = 467)) or
								((vState = 457) and (hState = 468)) or
								((vState = 457) and (hState = 469)) or
								((vState = 457) and (hState = 470)) or
								((vState = 457) and (hState = 471)) or
								((vState = 457) and (hState = 472)) or
								((vState = 457) and (hState = 473)) or
								((vState = 457) and (hState = 474)) or
								((vState = 457) and (hState = 475)) or
								((vState = 457) and (hState = 476)) or
								((vState = 457) and (hState = 477)) or
								((vState = 457) and (hState = 478)) or
								((vState = 457) and (hState = 479)) or
								((vState = 457) and (hState = 480)) or
								((vState = 457) and (hState = 481)) or
								((vState = 457) and (hState = 482)) or
								((vState = 457) and (hState = 511)) or
								((vState = 457) and (hState = 519)) or
								((vState = 457) and (hState = 520)) or
								((vState = 457) and (hState = 521)) or
								((vState = 457) and (hState = 522)) or
								((vState = 457) and (hState = 523)) or
								((vState = 457) and (hState = 524)) or
								((vState = 457) and (hState = 525)) or
								((vState = 457) and (hState = 526)) or
								((vState = 457) and (hState = 527)) or
								((vState = 457) and (hState = 531)) or
								((vState = 457) and (hState = 532)) or
								((vState = 457) and (hState = 533)) or
								((vState = 457) and (hState = 534)) or
								((vState = 457) and (hState = 574)) or
								((vState = 457) and (hState = 594)) or
								((vState = 457) and (hState = 595)) or
								((vState = 457) and (hState = 596)) or
								((vState = 458) and (hState = 287)) or
								((vState = 458) and (hState = 319)) or
								((vState = 458) and (hState = 334)) or
								((vState = 458) and (hState = 335)) or
								((vState = 458) and (hState = 336)) or
								((vState = 458) and (hState = 337)) or
								((vState = 458) and (hState = 338)) or
								((vState = 458) and (hState = 362)) or
								((vState = 458) and (hState = 384)) or
								((vState = 458) and (hState = 388)) or
								((vState = 458) and (hState = 418)) or
								((vState = 458) and (hState = 428)) or
								((vState = 458) and (hState = 439)) or
								((vState = 458) and (hState = 440)) or
								((vState = 458) and (hState = 441)) or
								((vState = 458) and (hState = 442)) or
								((vState = 458) and (hState = 443)) or
								((vState = 458) and (hState = 444)) or
								((vState = 458) and (hState = 445)) or
								((vState = 458) and (hState = 446)) or
								((vState = 458) and (hState = 447)) or
								((vState = 458) and (hState = 448)) or
								((vState = 458) and (hState = 449)) or
								((vState = 458) and (hState = 450)) or
								((vState = 458) and (hState = 451)) or
								((vState = 458) and (hState = 452)) or
								((vState = 458) and (hState = 453)) or
								((vState = 458) and (hState = 454)) or
								((vState = 458) and (hState = 455)) or
								((vState = 458) and (hState = 456)) or
								((vState = 458) and (hState = 457)) or
								((vState = 458) and (hState = 458)) or
								((vState = 458) and (hState = 459)) or
								((vState = 458) and (hState = 460)) or
								((vState = 458) and (hState = 461)) or
								((vState = 458) and (hState = 479)) or
								((vState = 458) and (hState = 480)) or
								((vState = 458) and (hState = 481)) or
								((vState = 458) and (hState = 482)) or
								((vState = 458) and (hState = 483)) or
								((vState = 458) and (hState = 484)) or
								((vState = 458) and (hState = 485)) or
								((vState = 458) and (hState = 486)) or
								((vState = 458) and (hState = 487)) or
								((vState = 458) and (hState = 492)) or
								((vState = 458) and (hState = 511)) or
								((vState = 458) and (hState = 512)) or
								((vState = 458) and (hState = 517)) or
								((vState = 458) and (hState = 518)) or
								((vState = 458) and (hState = 519)) or
								((vState = 458) and (hState = 520)) or
								((vState = 458) and (hState = 521)) or
								((vState = 458) and (hState = 522)) or
								((vState = 458) and (hState = 523)) or
								((vState = 458) and (hState = 531)) or
								((vState = 458) and (hState = 532)) or
								((vState = 458) and (hState = 533)) or
								((vState = 458) and (hState = 594)) or
								((vState = 459) and (hState = 319)) or
								((vState = 459) and (hState = 335)) or
								((vState = 459) and (hState = 336)) or
								((vState = 459) and (hState = 362)) or
								((vState = 459) and (hState = 384)) or
								((vState = 459) and (hState = 428)) or
								((vState = 459) and (hState = 449)) or
								((vState = 459) and (hState = 450)) or
								((vState = 459) and (hState = 459)) or
								((vState = 459) and (hState = 460)) or
								((vState = 459) and (hState = 479)) or
								((vState = 459) and (hState = 484)) or
								((vState = 459) and (hState = 485)) or
								((vState = 459) and (hState = 492)) or
								((vState = 459) and (hState = 511)) or
								((vState = 459) and (hState = 512)) or
								((vState = 459) and (hState = 521)) or
								((vState = 459) and (hState = 522)) or
								((vState = 459) and (hState = 531)) or
								((vState = 459) and (hState = 532)) or
								((vState = 459) and (hState = 594)) or
								((vState = 460) and (hState = 299)) or
								((vState = 460) and (hState = 300)) or
								((vState = 460) and (hState = 319)) or
								((vState = 460) and (hState = 335)) or
								((vState = 460) and (hState = 336)) or
								((vState = 460) and (hState = 362)) or
								((vState = 460) and (hState = 384)) or
								((vState = 460) and (hState = 392)) or
								((vState = 460) and (hState = 406)) or
								((vState = 460) and (hState = 428)) or
								((vState = 460) and (hState = 449)) or
								((vState = 460) and (hState = 459)) or
								((vState = 460) and (hState = 490)) or
								((vState = 460) and (hState = 511)) or
								((vState = 460) and (hState = 522)) or
								((vState = 460) and (hState = 594)) or
								((vState = 461) and (hState = 289)) or
								((vState = 461) and (hState = 299)) or
								((vState = 461) and (hState = 319)) or
								((vState = 461) and (hState = 335)) or
								((vState = 461) and (hState = 336)) or
								((vState = 461) and (hState = 354)) or
								((vState = 461) and (hState = 355)) or
								((vState = 461) and (hState = 362)) or
								((vState = 461) and (hState = 384)) or
								((vState = 461) and (hState = 385)) or
								((vState = 461) and (hState = 386)) or
								((vState = 461) and (hState = 387)) or
								((vState = 461) and (hState = 391)) or
								((vState = 461) and (hState = 402)) or
								((vState = 461) and (hState = 406)) or
								((vState = 461) and (hState = 416)) or
								((vState = 461) and (hState = 428)) or
								((vState = 461) and (hState = 437)) or
								((vState = 461) and (hState = 449)) or
								((vState = 461) and (hState = 459)) or
								((vState = 461) and (hState = 490)) or
								((vState = 461) and (hState = 496)) or
								((vState = 461) and (hState = 497)) or
								((vState = 461) and (hState = 511)) or
								((vState = 461) and (hState = 522)) or
								((vState = 461) and (hState = 530)) or
								((vState = 461) and (hState = 572)) or
								((vState = 461) and (hState = 585)) or
								((vState = 461) and (hState = 594)) or
								((vState = 462) and (hState = 299)) or
								((vState = 462) and (hState = 319)) or
								((vState = 462) and (hState = 335)) or
								((vState = 462) and (hState = 336)) or
								((vState = 462) and (hState = 341)) or
								((vState = 462) and (hState = 356)) or
								((vState = 462) and (hState = 357)) or
								((vState = 462) and (hState = 362)) or
								((vState = 462) and (hState = 371)) or
								((vState = 462) and (hState = 384)) or
								((vState = 462) and (hState = 385)) or
								((vState = 462) and (hState = 386)) or
								((vState = 462) and (hState = 387)) or
								((vState = 462) and (hState = 390)) or
								((vState = 462) and (hState = 404)) or
								((vState = 462) and (hState = 405)) or
								((vState = 462) and (hState = 406)) or
								((vState = 462) and (hState = 449)) or
								((vState = 462) and (hState = 458)) or
								((vState = 462) and (hState = 487)) or
								((vState = 462) and (hState = 488)) or
								((vState = 462) and (hState = 501)) or
								((vState = 462) and (hState = 502)) or
								((vState = 462) and (hState = 511)) or
								((vState = 462) and (hState = 522)) or
								((vState = 462) and (hState = 529)) or
								((vState = 462) and (hState = 530)) or
								((vState = 462) and (hState = 534)) or
								((vState = 462) and (hState = 584)) or
								((vState = 462) and (hState = 593)) or
								((vState = 463) and (hState = 299)) or
								((vState = 463) and (hState = 319)) or
								((vState = 463) and (hState = 335)) or
								((vState = 463) and (hState = 336)) or
								((vState = 463) and (hState = 337)) or
								((vState = 463) and (hState = 360)) or
								((vState = 463) and (hState = 361)) or
								((vState = 463) and (hState = 362)) or
								((vState = 463) and (hState = 384)) or
								((vState = 463) and (hState = 385)) or
								((vState = 463) and (hState = 390)) or
								((vState = 463) and (hState = 405)) or
								((vState = 463) and (hState = 406)) or
								((vState = 463) and (hState = 413)) or
								((vState = 463) and (hState = 427)) or
								((vState = 463) and (hState = 434)) or
								((vState = 463) and (hState = 448)) or
								((vState = 463) and (hState = 487)) or
								((vState = 463) and (hState = 488)) or
								((vState = 463) and (hState = 512)) or
								((vState = 463) and (hState = 515)) or
								((vState = 463) and (hState = 521)) or
								((vState = 463) and (hState = 522)) or
								((vState = 463) and (hState = 525)) or
								((vState = 463) and (hState = 526)) or
								((vState = 463) and (hState = 527)) or
								((vState = 463) and (hState = 528)) or
								((vState = 463) and (hState = 535)) or
								((vState = 463) and (hState = 536)) or
								((vState = 463) and (hState = 583)) or
								((vState = 463) and (hState = 593)) or
								((vState = 464) and (hState = 299)) or
								((vState = 464) and (hState = 319)) or
								((vState = 464) and (hState = 362)) or
								((vState = 464) and (hState = 384)) or
								((vState = 464) and (hState = 385)) or
								((vState = 464) and (hState = 427)) or
								((vState = 464) and (hState = 448)) or
								((vState = 464) and (hState = 512)) or
								((vState = 464) and (hState = 525)) or
								((vState = 464) and (hState = 536)) or
								((vState = 464) and (hState = 593)) or
								((vState = 465) and (hState = 319)) or
								((vState = 465) and (hState = 384)) or
								((vState = 465) and (hState = 407)) or
								((vState = 465) and (hState = 427)) or
								((vState = 465) and (hState = 455)) or
								((vState = 465) and (hState = 456)) or
								((vState = 465) and (hState = 476)) or
								((vState = 465) and (hState = 512)) or
								((vState = 465) and (hState = 593)) or
								((vState = 466) and (hState = 293)) or
								((vState = 466) and (hState = 298)) or
								((vState = 466) and (hState = 319)) or
								((vState = 466) and (hState = 334)) or
								((vState = 466) and (hState = 363)) or
								((vState = 466) and (hState = 364)) or
								((vState = 466) and (hState = 365)) or
								((vState = 466) and (hState = 366)) or
								((vState = 466) and (hState = 367)) or
								((vState = 466) and (hState = 368)) or
								((vState = 466) and (hState = 384)) or
								((vState = 466) and (hState = 388)) or
								((vState = 466) and (hState = 407)) or
								((vState = 466) and (hState = 408)) or
								((vState = 466) and (hState = 409)) or
								((vState = 466) and (hState = 410)) or
								((vState = 466) and (hState = 411)) or
								((vState = 466) and (hState = 427)) or
								((vState = 466) and (hState = 432)) or
								((vState = 466) and (hState = 454)) or
								((vState = 466) and (hState = 455)) or
								((vState = 466) and (hState = 456)) or
								((vState = 466) and (hState = 457)) or
								((vState = 466) and (hState = 458)) or
								((vState = 466) and (hState = 459)) or
								((vState = 466) and (hState = 460)) or
								((vState = 466) and (hState = 461)) or
								((vState = 466) and (hState = 462)) or
								((vState = 466) and (hState = 463)) or
								((vState = 466) and (hState = 464)) or
								((vState = 466) and (hState = 465)) or
								((vState = 466) and (hState = 466)) or
								((vState = 466) and (hState = 467)) or
								((vState = 466) and (hState = 476)) or
								((vState = 466) and (hState = 485)) or
								((vState = 466) and (hState = 491)) or
								((vState = 466) and (hState = 512)) or
								((vState = 466) and (hState = 517)) or
								((vState = 466) and (hState = 524)) or
								((vState = 466) and (hState = 537)) or
								((vState = 466) and (hState = 593)) or
								((vState = 467) and (hState = 294)) or
								((vState = 467) and (hState = 298)) or
								((vState = 467) and (hState = 319)) or
								((vState = 467) and (hState = 334)) or
								((vState = 467) and (hState = 340)) or
								((vState = 467) and (hState = 363)) or
								((vState = 467) and (hState = 367)) or
								((vState = 467) and (hState = 368)) or
								((vState = 467) and (hState = 384)) or
								((vState = 467) and (hState = 388)) or
								((vState = 467) and (hState = 407)) or
								((vState = 467) and (hState = 408)) or
								((vState = 467) and (hState = 409)) or
								((vState = 467) and (hState = 410)) or
								((vState = 467) and (hState = 411)) or
								((vState = 467) and (hState = 427)) or
								((vState = 467) and (hState = 453)) or
								((vState = 467) and (hState = 458)) or
								((vState = 467) and (hState = 469)) or
								((vState = 467) and (hState = 470)) or
								((vState = 467) and (hState = 475)) or
								((vState = 467) and (hState = 492)) or
								((vState = 467) and (hState = 518)) or
								((vState = 467) and (hState = 519)) or
								((vState = 467) and (hState = 520)) or
								((vState = 467) and (hState = 521)) or
								((vState = 467) and (hState = 522)) or
								((vState = 467) and (hState = 523)) or
								((vState = 467) and (hState = 568)) or
								((vState = 468) and (hState = 298)) or
								((vState = 468) and (hState = 345)) or
								((vState = 468) and (hState = 363)) or
								((vState = 468) and (hState = 367)) or
								((vState = 468) and (hState = 368)) or
								((vState = 468) and (hState = 369)) or
								((vState = 468) and (hState = 370)) or
								((vState = 468) and (hState = 371)) or
								((vState = 468) and (hState = 383)) or
								((vState = 468) and (hState = 384)) or
								((vState = 468) and (hState = 385)) or
								((vState = 468) and (hState = 386)) or
								((vState = 468) and (hState = 387)) or
								((vState = 468) and (hState = 407)) or
								((vState = 468) and (hState = 408)) or
								((vState = 468) and (hState = 409)) or
								((vState = 468) and (hState = 410)) or
								((vState = 468) and (hState = 411)) or
								((vState = 468) and (hState = 427)) or
								((vState = 468) and (hState = 428)) or
								((vState = 468) and (hState = 429)) or
								((vState = 468) and (hState = 473)) or
								((vState = 468) and (hState = 474)) or
								((vState = 468) and (hState = 475)) or
								((vState = 468) and (hState = 513)) or
								((vState = 468) and (hState = 519)) or
								((vState = 468) and (hState = 520)) or
								((vState = 468) and (hState = 567)) or
								((vState = 468) and (hState = 579)) or
								((vState = 469) and (hState = 298)) or
								((vState = 469) and (hState = 345)) or
								((vState = 469) and (hState = 363)) or
								((vState = 469) and (hState = 383)) or
								((vState = 469) and (hState = 384)) or
								((vState = 469) and (hState = 385)) or
								((vState = 469) and (hState = 407)) or
								((vState = 469) and (hState = 408)) or
								((vState = 469) and (hState = 409)) or
								((vState = 469) and (hState = 427)) or
								((vState = 469) and (hState = 428)) or
								((vState = 469) and (hState = 474)) or
								((vState = 469) and (hState = 475)) or
								((vState = 469) and (hState = 513)) or
								((vState = 469) and (hState = 519)) or
								((vState = 469) and (hState = 520)) or
								((vState = 470) and (hState = 297)) or
								((vState = 470) and (hState = 298)) or
								((vState = 470) and (hState = 345)) or
								((vState = 470) and (hState = 363)) or
								((vState = 470) and (hState = 364)) or
								((vState = 470) and (hState = 383)) or
								((vState = 470) and (hState = 384)) or
								((vState = 470) and (hState = 408)) or
								((vState = 470) and (hState = 426)) or
								((vState = 470) and (hState = 427)) or
								((vState = 470) and (hState = 445)) or
								((vState = 470) and (hState = 474)) or
								((vState = 470) and (hState = 481)) or
								((vState = 470) and (hState = 513)) or
								((vState = 470) and (hState = 519)) or
								((vState = 470) and (hState = 520)) or
								((vState = 471) and (hState = 297)) or
								((vState = 471) and (hState = 298)) or
								((vState = 471) and (hState = 343)) or
								((vState = 471) and (hState = 344)) or
								((vState = 471) and (hState = 345)) or
								((vState = 471) and (hState = 346)) or
								((vState = 471) and (hState = 363)) or
								((vState = 471) and (hState = 364)) or
								((vState = 471) and (hState = 381)) or
								((vState = 471) and (hState = 382)) or
								((vState = 471) and (hState = 383)) or
								((vState = 471) and (hState = 384)) or
								((vState = 471) and (hState = 426)) or
								((vState = 471) and (hState = 427)) or
								((vState = 471) and (hState = 444)) or
								((vState = 471) and (hState = 445)) or
								((vState = 471) and (hState = 460)) or
								((vState = 471) and (hState = 474)) or
								((vState = 471) and (hState = 478)) or
								((vState = 471) and (hState = 479)) or
								((vState = 471) and (hState = 480)) or
								((vState = 471) and (hState = 481)) or
								((vState = 471) and (hState = 513)) or
								((vState = 471) and (hState = 518)) or
								((vState = 471) and (hState = 519)) or
								((vState = 471) and (hState = 520)) or
								((vState = 471) and (hState = 541)) or
								((vState = 472) and (hState = 298)) or
								((vState = 472) and (hState = 325)) or
								((vState = 472) and (hState = 326)) or
								((vState = 472) and (hState = 331)) or
								((vState = 472) and (hState = 332)) or
								((vState = 472) and (hState = 333)) or
								((vState = 472) and (hState = 334)) or
								((vState = 472) and (hState = 363)) or
								((vState = 472) and (hState = 364)) or
								((vState = 472) and (hState = 378)) or
								((vState = 472) and (hState = 379)) or
								((vState = 472) and (hState = 380)) or
								((vState = 472) and (hState = 381)) or
								((vState = 472) and (hState = 382)) or
								((vState = 472) and (hState = 383)) or
								((vState = 472) and (hState = 384)) or
								((vState = 472) and (hState = 416)) or
								((vState = 472) and (hState = 444)) or
								((vState = 472) and (hState = 445)) or
								((vState = 472) and (hState = 446)) or
								((vState = 472) and (hState = 481)) or
								((vState = 472) and (hState = 482)) or
								((vState = 472) and (hState = 514)) or
								((vState = 472) and (hState = 515)) or
								((vState = 472) and (hState = 519)) or
								((vState = 472) and (hState = 520)) or
								((vState = 472) and (hState = 521)) or
								((vState = 472) and (hState = 522)) or
								((vState = 473) and (hState = 299)) or
								((vState = 473) and (hState = 329)) or
								((vState = 473) and (hState = 330)) or
								((vState = 473) and (hState = 331)) or
								((vState = 473) and (hState = 332)) or
								((vState = 473) and (hState = 333)) or
								((vState = 473) and (hState = 334)) or
								((vState = 473) and (hState = 335)) or
								((vState = 473) and (hState = 336)) or
								((vState = 473) and (hState = 337)) or
								((vState = 473) and (hState = 347)) or
								((vState = 473) and (hState = 380)) or
								((vState = 473) and (hState = 381)) or
								((vState = 473) and (hState = 382)) or
								((vState = 473) and (hState = 383)) or
								((vState = 473) and (hState = 384)) or
								((vState = 473) and (hState = 402)) or
								((vState = 473) and (hState = 417)) or
								((vState = 473) and (hState = 443)) or
								((vState = 473) and (hState = 444)) or
								((vState = 473) and (hState = 445)) or
								((vState = 473) and (hState = 484)) or
								((vState = 473) and (hState = 485)) or
								((vState = 473) and (hState = 486)) or
								((vState = 473) and (hState = 487)) or
								((vState = 473) and (hState = 523)) or
								((vState = 473) and (hState = 542)) or
								((vState = 473) and (hState = 562)) or
								((vState = 473) and (hState = 563)) or
								((vState = 473) and (hState = 564)) or
								((vState = 473) and (hState = 590)) or
								((vState = 474) and (hState = 333)) or
								((vState = 474) and (hState = 334)) or
								((vState = 474) and (hState = 335)) or
								((vState = 474) and (hState = 336)) or
								((vState = 474) and (hState = 337)) or
								((vState = 474) and (hState = 347)) or
								((vState = 474) and (hState = 381)) or
								((vState = 474) and (hState = 382)) or
								((vState = 474) and (hState = 383)) or
								((vState = 474) and (hState = 384)) or
								((vState = 474) and (hState = 426)) or
								((vState = 474) and (hState = 443)) or
								((vState = 474) and (hState = 444)) or
								((vState = 474) and (hState = 472)) or
								((vState = 474) and (hState = 473)) or
								((vState = 474) and (hState = 514)) or
								((vState = 474) and (hState = 562)) or
								((vState = 474) and (hState = 563)) or
								((vState = 474) and (hState = 564)) or
								((vState = 474) and (hState = 590)) or
								((vState = 475) and (hState = 336)) or
								((vState = 475) and (hState = 337)) or
								((vState = 475) and (hState = 338)) or
								((vState = 475) and (hState = 339)) or
								((vState = 475) and (hState = 340)) or
								((vState = 475) and (hState = 345)) or
								((vState = 475) and (hState = 346)) or
								((vState = 475) and (hState = 347)) or
								((vState = 475) and (hState = 348)) or
								((vState = 475) and (hState = 381)) or
								((vState = 475) and (hState = 382)) or
								((vState = 475) and (hState = 383)) or
								((vState = 475) and (hState = 442)) or
								((vState = 475) and (hState = 443)) or
								((vState = 475) and (hState = 471)) or
								((vState = 475) and (hState = 472)) or
								((vState = 475) and (hState = 473)) or
								((vState = 475) and (hState = 474)) or
								((vState = 475) and (hState = 501)) or
								((vState = 475) and (hState = 514)) or
								((vState = 475) and (hState = 518)) or
								((vState = 475) and (hState = 562)) or
								((vState = 475) and (hState = 590)) or
								((vState = 476) and (hState = 339)) or
								((vState = 476) and (hState = 340)) or
								((vState = 476) and (hState = 341)) or
								((vState = 476) and (hState = 342)) or
								((vState = 476) and (hState = 343)) or
								((vState = 476) and (hState = 344)) or
								((vState = 476) and (hState = 345)) or
								((vState = 476) and (hState = 346)) or
								((vState = 476) and (hState = 347)) or
								((vState = 476) and (hState = 348)) or
								((vState = 476) and (hState = 380)) or
								((vState = 476) and (hState = 381)) or
								((vState = 476) and (hState = 382)) or
								((vState = 476) and (hState = 383)) or
								((vState = 476) and (hState = 421)) or
								((vState = 476) and (hState = 422)) or
								((vState = 476) and (hState = 442)) or
								((vState = 476) and (hState = 471)) or
								((vState = 476) and (hState = 472)) or
								((vState = 476) and (hState = 473)) or
								((vState = 476) and (hState = 501)) or
								((vState = 476) and (hState = 502)) or
								((vState = 476) and (hState = 518)) or
								((vState = 477) and (hState = 340)) or
								((vState = 477) and (hState = 341)) or
								((vState = 477) and (hState = 342)) or
								((vState = 477) and (hState = 343)) or
								((vState = 477) and (hState = 344)) or
								((vState = 477) and (hState = 345)) or
								((vState = 477) and (hState = 346)) or
								((vState = 477) and (hState = 347)) or
								((vState = 477) and (hState = 348)) or
								((vState = 477) and (hState = 349)) or
								((vState = 477) and (hState = 350)) or
								((vState = 477) and (hState = 379)) or
								((vState = 477) and (hState = 380)) or
								((vState = 477) and (hState = 381)) or
								((vState = 477) and (hState = 382)) or
								((vState = 477) and (hState = 383)) or
								((vState = 477) and (hState = 389)) or
								((vState = 477) and (hState = 421)) or
								((vState = 477) and (hState = 422)) or
								((vState = 477) and (hState = 470)) or
								((vState = 477) and (hState = 471)) or
								((vState = 477) and (hState = 472)) or
								((vState = 477) and (hState = 500)) or
								((vState = 477) and (hState = 501)) or
								((vState = 477) and (hState = 502)) or
								((vState = 477) and (hState = 503)) or
								((vState = 477) and (hState = 518)) or
								((vState = 477) and (hState = 525)) or
								((vState = 477) and (hState = 556)) or
								((vState = 477) and (hState = 572)) or
								((vState = 478) and (hState = 303)) or
								((vState = 478) and (hState = 344)) or
								((vState = 478) and (hState = 345)) or
								((vState = 478) and (hState = 346)) or
								((vState = 478) and (hState = 347)) or
								((vState = 478) and (hState = 348)) or
								((vState = 478) and (hState = 349)) or
								((vState = 478) and (hState = 350)) or
								((vState = 478) and (hState = 379)) or
								((vState = 478) and (hState = 383)) or
								((vState = 478) and (hState = 391)) or
								((vState = 478) and (hState = 397)) or
								((vState = 478) and (hState = 421)) or
								((vState = 478) and (hState = 422)) or
								((vState = 478) and (hState = 423)) or
								((vState = 478) and (hState = 466)) or
								((vState = 478) and (hState = 470)) or
								((vState = 478) and (hState = 471)) or
								((vState = 478) and (hState = 505)) or
								((vState = 478) and (hState = 506)) or
								((vState = 478) and (hState = 507)) or
								((vState = 478) and (hState = 516)) or
								((vState = 478) and (hState = 517)) or
								((vState = 478) and (hState = 526)) or
								((vState = 478) and (hState = 527)) or
								((vState = 478) and (hState = 553)) or
								((vState = 478) and (hState = 585)) or
								((vState = 478) and (hState = 589)) or
								((vState = 479) and (hState = 347)) or
								((vState = 479) and (hState = 348)) or
								((vState = 479) and (hState = 349)) or
								((vState = 479) and (hState = 350)) or
								((vState = 479) and (hState = 351)) or
								((vState = 479) and (hState = 352)) or
								((vState = 479) and (hState = 378)) or
								((vState = 479) and (hState = 379)) or
								((vState = 479) and (hState = 383)) or
								((vState = 479) and (hState = 394)) or
								((vState = 479) and (hState = 395)) or
								((vState = 479) and (hState = 396)) or
								((vState = 479) and (hState = 439)) or
								((vState = 479) and (hState = 468)) or
								((vState = 479) and (hState = 469)) or
								((vState = 479) and (hState = 470)) or
								((vState = 479) and (hState = 505)) or
								((vState = 479) and (hState = 506)) or
								((vState = 479) and (hState = 516)) or
								((vState = 479) and (hState = 517)) or
								((vState = 479) and (hState = 552)) or
								((vState = 479) and (hState = 569)) or
								((vState = 479) and (hState = 585)) or
								((vState = 479) and (hState = 589)) or
								((vState = 480) and (hState = 350)) or
								((vState = 480) and (hState = 351)) or
								((vState = 480) and (hState = 352)) or
								((vState = 480) and (hState = 378)) or
								((vState = 480) and (hState = 383)) or
								((vState = 480) and (hState = 468)) or
								((vState = 480) and (hState = 469)) or
								((vState = 480) and (hState = 470)) or
								((vState = 480) and (hState = 504)) or
								((vState = 480) and (hState = 516)) or
								((vState = 480) and (hState = 517)) or
								((vState = 480) and (hState = 585)) or
								((vState = 480) and (hState = 589)) or
								((vState = 481) and (hState = 350)) or
								((vState = 481) and (hState = 351)) or
								((vState = 481) and (hState = 352)) or
								((vState = 481) and (hState = 353)) or
								((vState = 481) and (hState = 354)) or
								((vState = 481) and (hState = 355)) or
								((vState = 481) and (hState = 383)) or
								((vState = 481) and (hState = 469)) or
								((vState = 481) and (hState = 470)) or
								((vState = 481) and (hState = 516)) or
								((vState = 481) and (hState = 517)) or
								((vState = 481) and (hState = 528)) or
								((vState = 481) and (hState = 542)) or
								((vState = 481) and (hState = 584)) or
								((vState = 481) and (hState = 585)) or
								((vState = 482) and (hState = 350)) or
								((vState = 482) and (hState = 351)) or
								((vState = 482) and (hState = 352)) or
								((vState = 482) and (hState = 353)) or
								((vState = 482) and (hState = 354)) or
								((vState = 482) and (hState = 355)) or
								((vState = 482) and (hState = 356)) or
								((vState = 482) and (hState = 357)) or
								((vState = 482) and (hState = 358)) or
								((vState = 482) and (hState = 376)) or
								((vState = 482) and (hState = 377)) or
								((vState = 482) and (hState = 383)) or
								((vState = 482) and (hState = 409)) or
								((vState = 482) and (hState = 417)) or
								((vState = 482) and (hState = 428)) or
								((vState = 482) and (hState = 437)) or
								((vState = 482) and (hState = 469)) or
								((vState = 482) and (hState = 470)) or
								((vState = 482) and (hState = 502)) or
								((vState = 482) and (hState = 516)) or
								((vState = 482) and (hState = 517)) or
								((vState = 482) and (hState = 528)) or
								((vState = 482) and (hState = 542)) or
								((vState = 482) and (hState = 547)) or
								((vState = 482) and (hState = 548)) or
								((vState = 482) and (hState = 558)) or
								((vState = 482) and (hState = 584)) or
								((vState = 482) and (hState = 585)) or
								((vState = 483) and (hState = 344)) or
								((vState = 483) and (hState = 345)) or
								((vState = 483) and (hState = 346)) or
								((vState = 483) and (hState = 347)) or
								((vState = 483) and (hState = 348)) or
								((vState = 483) and (hState = 349)) or
								((vState = 483) and (hState = 350)) or
								((vState = 483) and (hState = 359)) or
								((vState = 483) and (hState = 360)) or
								((vState = 483) and (hState = 361)) or
								((vState = 483) and (hState = 373)) or
								((vState = 483) and (hState = 374)) or
								((vState = 483) and (hState = 375)) or
								((vState = 483) and (hState = 383)) or
								((vState = 483) and (hState = 406)) or
								((vState = 483) and (hState = 407)) or
								((vState = 483) and (hState = 416)) or
								((vState = 483) and (hState = 429)) or
								((vState = 483) and (hState = 471)) or
								((vState = 483) and (hState = 501)) or
								((vState = 483) and (hState = 525)) or
								((vState = 483) and (hState = 542)) or
								((vState = 483) and (hState = 546)) or
								((vState = 483) and (hState = 557)) or
								((vState = 483) and (hState = 566)) or
								((vState = 483) and (hState = 567)) or
								((vState = 483) and (hState = 583)) or
								((vState = 483) and (hState = 584)) or
								((vState = 483) and (hState = 585)) or
								((vState = 483) and (hState = 586)) or
								((vState = 483) and (hState = 587)) or
								((vState = 483) and (hState = 588)) or
								((vState = 484) and (hState = 308)) or
								((vState = 484) and (hState = 315)) or
								((vState = 484) and (hState = 316)) or
								((vState = 484) and (hState = 317)) or
								((vState = 484) and (hState = 318)) or
								((vState = 484) and (hState = 319)) or
								((vState = 484) and (hState = 320)) or
								((vState = 484) and (hState = 321)) or
								((vState = 484) and (hState = 322)) or
								((vState = 484) and (hState = 323)) or
								((vState = 484) and (hState = 324)) or
								((vState = 484) and (hState = 325)) or
								((vState = 484) and (hState = 326)) or
								((vState = 484) and (hState = 327)) or
								((vState = 484) and (hState = 328)) or
								((vState = 484) and (hState = 329)) or
								((vState = 484) and (hState = 330)) or
								((vState = 484) and (hState = 331)) or
								((vState = 484) and (hState = 335)) or
								((vState = 484) and (hState = 336)) or
								((vState = 484) and (hState = 337)) or
								((vState = 484) and (hState = 338)) or
								((vState = 484) and (hState = 339)) or
								((vState = 484) and (hState = 340)) or
								((vState = 484) and (hState = 362)) or
								((vState = 484) and (hState = 363)) or
								((vState = 484) and (hState = 364)) or
								((vState = 484) and (hState = 372)) or
								((vState = 484) and (hState = 375)) or
								((vState = 484) and (hState = 383)) or
								((vState = 484) and (hState = 404)) or
								((vState = 484) and (hState = 405)) or
								((vState = 484) and (hState = 431)) or
								((vState = 484) and (hState = 432)) or
								((vState = 484) and (hState = 433)) or
								((vState = 484) and (hState = 524)) or
								((vState = 484) and (hState = 542)) or
								((vState = 484) and (hState = 543)) or
								((vState = 484) and (hState = 557)) or
								((vState = 484) and (hState = 583)) or
								((vState = 484) and (hState = 584)) or
								((vState = 484) and (hState = 588)) or
								((vState = 485) and (hState = 317)) or
								((vState = 485) and (hState = 318)) or
								((vState = 485) and (hState = 383)) or
								((vState = 485) and (hState = 431)) or
								((vState = 485) and (hState = 432)) or
								((vState = 485) and (hState = 433)) or
								((vState = 485) and (hState = 542)) or
								((vState = 485) and (hState = 557)) or
								((vState = 485) and (hState = 583)) or
								((vState = 485) and (hState = 584)) or
								((vState = 485) and (hState = 588)) or
								((vState = 486) and (hState = 318)) or
								((vState = 486) and (hState = 383)) or
								((vState = 486) and (hState = 431)) or
								((vState = 486) and (hState = 541)) or
								((vState = 486) and (hState = 542)) or
								((vState = 486) and (hState = 556)) or
								((vState = 486) and (hState = 557)) or
								((vState = 486) and (hState = 584)) or
								((vState = 487) and (hState = 309)) or
								((vState = 487) and (hState = 318)) or
								((vState = 487) and (hState = 356)) or
								((vState = 487) and (hState = 368)) or
								((vState = 487) and (hState = 383)) or
								((vState = 487) and (hState = 400)) or
								((vState = 487) and (hState = 412)) or
								((vState = 487) and (hState = 434)) or
								((vState = 487) and (hState = 474)) or
								((vState = 487) and (hState = 485)) or
								((vState = 487) and (hState = 486)) or
								((vState = 487) and (hState = 487)) or
								((vState = 487) and (hState = 496)) or
								((vState = 487) and (hState = 520)) or
								((vState = 487) and (hState = 540)) or
								((vState = 487) and (hState = 541)) or
								((vState = 487) and (hState = 542)) or
								((vState = 487) and (hState = 555)) or
								((vState = 487) and (hState = 556)) or
								((vState = 487) and (hState = 557)) or
								((vState = 487) and (hState = 558)) or
								((vState = 487) and (hState = 559)) or
								((vState = 487) and (hState = 560)) or
								((vState = 487) and (hState = 561)) or
								((vState = 487) and (hState = 562)) or
								((vState = 487) and (hState = 563)) or
								((vState = 487) and (hState = 564)) or
								((vState = 487) and (hState = 584)) or
								((vState = 488) and (hState = 310)) or
								((vState = 488) and (hState = 319)) or
								((vState = 488) and (hState = 366)) or
								((vState = 488) and (hState = 383)) or
								((vState = 488) and (hState = 397)) or
								((vState = 488) and (hState = 411)) or
								((vState = 488) and (hState = 429)) or
								((vState = 488) and (hState = 430)) or
								((vState = 488) and (hState = 434)) or
								((vState = 488) and (hState = 435)) or
								((vState = 488) and (hState = 475)) or
								((vState = 488) and (hState = 489)) or
								((vState = 488) and (hState = 490)) or
								((vState = 488) and (hState = 491)) or
								((vState = 488) and (hState = 492)) or
								((vState = 488) and (hState = 493)) or
								((vState = 488) and (hState = 494)) or
								((vState = 488) and (hState = 518)) or
								((vState = 488) and (hState = 519)) or
								((vState = 488) and (hState = 520)) or
								((vState = 488) and (hState = 534)) or
								((vState = 488) and (hState = 535)) or
								((vState = 488) and (hState = 536)) or
								((vState = 488) and (hState = 537)) or
								((vState = 488) and (hState = 538)) or
								((vState = 488) and (hState = 539)) or
								((vState = 488) and (hState = 540)) or
								((vState = 488) and (hState = 541)) or
								((vState = 488) and (hState = 542)) or
								((vState = 488) and (hState = 543)) or
								((vState = 488) and (hState = 544)) or
								((vState = 488) and (hState = 545)) or
								((vState = 488) and (hState = 546)) or
								((vState = 488) and (hState = 547)) or
								((vState = 488) and (hState = 548)) or
								((vState = 488) and (hState = 549)) or
								((vState = 488) and (hState = 550)) or
								((vState = 488) and (hState = 551)) or
								((vState = 488) and (hState = 552)) or
								((vState = 488) and (hState = 553)) or
								((vState = 488) and (hState = 554)) or
								((vState = 488) and (hState = 584)) or
								((vState = 488) and (hState = 585)) or
								((vState = 488) and (hState = 586)) or
								((vState = 489) and (hState = 320)) or
								((vState = 489) and (hState = 357)) or
								((vState = 489) and (hState = 363)) or
								((vState = 489) and (hState = 373)) or
								((vState = 489) and (hState = 383)) or
								((vState = 489) and (hState = 395)) or
								((vState = 489) and (hState = 429)) or
								((vState = 489) and (hState = 430)) or
								((vState = 489) and (hState = 431)) or
								((vState = 489) and (hState = 432)) or
								((vState = 489) and (hState = 433)) or
								((vState = 489) and (hState = 434)) or
								((vState = 489) and (hState = 435)) or
								((vState = 489) and (hState = 436)) or
								((vState = 489) and (hState = 437)) or
								((vState = 489) and (hState = 476)) or
								((vState = 489) and (hState = 490)) or
								((vState = 489) and (hState = 491)) or
								((vState = 489) and (hState = 492)) or
								((vState = 489) and (hState = 493)) or
								((vState = 489) and (hState = 494)) or
								((vState = 489) and (hState = 517)) or
								((vState = 489) and (hState = 518)) or
								((vState = 489) and (hState = 519)) or
								((vState = 489) and (hState = 520)) or
								((vState = 489) and (hState = 521)) or
								((vState = 489) and (hState = 522)) or
								((vState = 489) and (hState = 523)) or
								((vState = 489) and (hState = 524)) or
								((vState = 489) and (hState = 525)) or
								((vState = 489) and (hState = 526)) or
								((vState = 489) and (hState = 527)) or
								((vState = 489) and (hState = 528)) or
								((vState = 489) and (hState = 529)) or
								((vState = 489) and (hState = 530)) or
								((vState = 489) and (hState = 534)) or
								((vState = 489) and (hState = 535)) or
								((vState = 489) and (hState = 536)) or
								((vState = 489) and (hState = 537)) or
								((vState = 489) and (hState = 538)) or
								((vState = 489) and (hState = 539)) or
								((vState = 489) and (hState = 540)) or
								((vState = 489) and (hState = 541)) or
								((vState = 489) and (hState = 542)) or
								((vState = 489) and (hState = 543)) or
								((vState = 489) and (hState = 544)) or
								((vState = 489) and (hState = 545)) or
								((vState = 489) and (hState = 546)) or
								((vState = 489) and (hState = 547)) or
								((vState = 489) and (hState = 552)) or
								((vState = 489) and (hState = 553)) or
								((vState = 489) and (hState = 554)) or
								((vState = 489) and (hState = 584)) or
								((vState = 489) and (hState = 585)) or
								((vState = 489) and (hState = 586)) or
								((vState = 490) and (hState = 383)) or
								((vState = 490) and (hState = 437)) or
								((vState = 490) and (hState = 490)) or
								((vState = 490) and (hState = 495)) or
								((vState = 490) and (hState = 526)) or
								((vState = 490) and (hState = 527)) or
								((vState = 490) and (hState = 528)) or
								((vState = 490) and (hState = 529)) or
								((vState = 490) and (hState = 530)) or
								((vState = 490) and (hState = 534)) or
								((vState = 490) and (hState = 535)) or
								((vState = 490) and (hState = 536)) or
								((vState = 490) and (hState = 537)) or
								((vState = 490) and (hState = 538)) or
								((vState = 490) and (hState = 539)) or
								((vState = 490) and (hState = 540)) or
								((vState = 490) and (hState = 552)) or
								((vState = 490) and (hState = 584)) or
								((vState = 490) and (hState = 585)) or
								((vState = 490) and (hState = 586)) or
								((vState = 491) and (hState = 383)) or
								((vState = 491) and (hState = 440)) or
								((vState = 491) and (hState = 500)) or
								((vState = 491) and (hState = 501)) or
								((vState = 491) and (hState = 502)) or
								((vState = 491) and (hState = 503)) or
								((vState = 491) and (hState = 504)) or
								((vState = 491) and (hState = 505)) or
								((vState = 491) and (hState = 506)) or
								((vState = 491) and (hState = 510)) or
								((vState = 491) and (hState = 511)) or
								((vState = 491) and (hState = 512)) or
								((vState = 491) and (hState = 513)) or
								((vState = 491) and (hState = 527)) or
								((vState = 491) and (hState = 528)) or
								((vState = 491) and (hState = 529)) or
								((vState = 491) and (hState = 530)) or
								((vState = 491) and (hState = 540)) or
								((vState = 491) and (hState = 552)) or
								((vState = 491) and (hState = 584)) or
								((vState = 491) and (hState = 585)) or
								((vState = 492) and (hState = 358)) or
								((vState = 492) and (hState = 359)) or
								((vState = 492) and (hState = 372)) or
								((vState = 492) and (hState = 407)) or
								((vState = 492) and (hState = 441)) or
								((vState = 492) and (hState = 442)) or
								((vState = 492) and (hState = 443)) or
								((vState = 492) and (hState = 444)) or
								((vState = 492) and (hState = 445)) or
								((vState = 492) and (hState = 502)) or
								((vState = 492) and (hState = 503)) or
								((vState = 492) and (hState = 504)) or
								((vState = 492) and (hState = 505)) or
								((vState = 492) and (hState = 506)) or
								((vState = 492) and (hState = 511)) or
								((vState = 492) and (hState = 512)) or
								((vState = 492) and (hState = 513)) or
								((vState = 492) and (hState = 527)) or
								((vState = 492) and (hState = 528)) or
								((vState = 492) and (hState = 529)) or
								((vState = 492) and (hState = 530)) or
								((vState = 492) and (hState = 531)) or
								((vState = 492) and (hState = 552)) or
								((vState = 492) and (hState = 584)) or
								((vState = 492) and (hState = 585)) or
								((vState = 493) and (hState = 314)) or
								((vState = 493) and (hState = 357)) or
								((vState = 493) and (hState = 358)) or
								((vState = 493) and (hState = 359)) or
								((vState = 493) and (hState = 372)) or
								((vState = 493) and (hState = 388)) or
								((vState = 493) and (hState = 406)) or
								((vState = 493) and (hState = 442)) or
								((vState = 493) and (hState = 443)) or
								((vState = 493) and (hState = 444)) or
								((vState = 493) and (hState = 449)) or
								((vState = 493) and (hState = 450)) or
								((vState = 493) and (hState = 451)) or
								((vState = 493) and (hState = 452)) or
								((vState = 493) and (hState = 453)) or
								((vState = 493) and (hState = 487)) or
								((vState = 493) and (hState = 503)) or
								((vState = 493) and (hState = 504)) or
								((vState = 493) and (hState = 505)) or
								((vState = 493) and (hState = 506)) or
								((vState = 493) and (hState = 511)) or
								((vState = 493) and (hState = 512)) or
								((vState = 493) and (hState = 513)) or
								((vState = 493) and (hState = 519)) or
								((vState = 493) and (hState = 520)) or
								((vState = 493) and (hState = 521)) or
								((vState = 493) and (hState = 522)) or
								((vState = 493) and (hState = 523)) or
								((vState = 493) and (hState = 524)) or
								((vState = 493) and (hState = 528)) or
								((vState = 493) and (hState = 529)) or
								((vState = 493) and (hState = 530)) or
								((vState = 493) and (hState = 551)) or
								((vState = 493) and (hState = 562)) or
								((vState = 493) and (hState = 578)) or
								((vState = 493) and (hState = 584)) or
								((vState = 493) and (hState = 585)) or
								((vState = 494) and (hState = 315)) or
								((vState = 494) and (hState = 356)) or
								((vState = 494) and (hState = 371)) or
								((vState = 494) and (hState = 385)) or
								((vState = 494) and (hState = 386)) or
								((vState = 494) and (hState = 387)) or
								((vState = 494) and (hState = 388)) or
								((vState = 494) and (hState = 405)) or
								((vState = 494) and (hState = 443)) or
								((vState = 494) and (hState = 444)) or
								((vState = 494) and (hState = 455)) or
								((vState = 494) and (hState = 456)) or
								((vState = 494) and (hState = 457)) or
								((vState = 494) and (hState = 458)) or
								((vState = 494) and (hState = 459)) or
								((vState = 494) and (hState = 480)) or
								((vState = 494) and (hState = 485)) or
								((vState = 494) and (hState = 507)) or
								((vState = 494) and (hState = 508)) or
								((vState = 494) and (hState = 509)) or
								((vState = 494) and (hState = 510)) or
								((vState = 494) and (hState = 511)) or
								((vState = 494) and (hState = 512)) or
								((vState = 494) and (hState = 513)) or
								((vState = 494) and (hState = 514)) or
								((vState = 494) and (hState = 515)) or
								((vState = 494) and (hState = 516)) or
								((vState = 494) and (hState = 517)) or
								((vState = 494) and (hState = 528)) or
								((vState = 494) and (hState = 577)) or
								((vState = 494) and (hState = 583)) or
								((vState = 494) and (hState = 584)) or
								((vState = 494) and (hState = 585)) or
								((vState = 494) and (hState = 595)) or
								((vState = 495) and (hState = 371)) or
								((vState = 495) and (hState = 385)) or
								((vState = 495) and (hState = 386)) or
								((vState = 495) and (hState = 387)) or
								((vState = 495) and (hState = 388)) or
								((vState = 495) and (hState = 507)) or
								((vState = 495) and (hState = 508)) or
								((vState = 495) and (hState = 509)) or
								((vState = 495) and (hState = 577)) or
								((vState = 495) and (hState = 583)) or
								((vState = 495) and (hState = 584)) or
								((vState = 495) and (hState = 585)) or
								((vState = 496) and (hState = 371)) or
								((vState = 496) and (hState = 383)) or
								((vState = 496) and (hState = 384)) or
								((vState = 496) and (hState = 390)) or
								((vState = 496) and (hState = 391)) or
								((vState = 496) and (hState = 392)) or
								((vState = 496) and (hState = 481)) or
								((vState = 496) and (hState = 482)) or
								((vState = 496) and (hState = 483)) or
								((vState = 496) and (hState = 577)) or
								((vState = 496) and (hState = 583)) or
								((vState = 496) and (hState = 584)) or
								((vState = 496) and (hState = 585)) or
								((vState = 496) and (hState = 594)) or
								((vState = 497) and (hState = 370)) or
								((vState = 497) and (hState = 371)) or
								((vState = 497) and (hState = 382)) or
								((vState = 497) and (hState = 383)) or
								((vState = 497) and (hState = 390)) or
								((vState = 497) and (hState = 483)) or
								((vState = 497) and (hState = 536)) or
								((vState = 497) and (hState = 537)) or
								((vState = 497) and (hState = 538)) or
								((vState = 497) and (hState = 539)) or
								((vState = 497) and (hState = 548)) or
								((vState = 497) and (hState = 569)) or
								((vState = 497) and (hState = 576)) or
								((vState = 497) and (hState = 577)) or
								((vState = 497) and (hState = 583)) or
								((vState = 497) and (hState = 584)) or
								((vState = 497) and (hState = 585)) or
								((vState = 497) and (hState = 594)) or
								((vState = 498) and (hState = 330)) or
								((vState = 498) and (hState = 350)) or
								((vState = 498) and (hState = 370)) or
								((vState = 498) and (hState = 371)) or
								((vState = 498) and (hState = 372)) or
								((vState = 498) and (hState = 373)) or
								((vState = 498) and (hState = 374)) or
								((vState = 498) and (hState = 375)) or
								((vState = 498) and (hState = 376)) or
								((vState = 498) and (hState = 377)) or
								((vState = 498) and (hState = 378)) or
								((vState = 498) and (hState = 383)) or
								((vState = 498) and (hState = 390)) or
								((vState = 498) and (hState = 401)) or
								((vState = 498) and (hState = 450)) or
								((vState = 498) and (hState = 474)) or
								((vState = 498) and (hState = 475)) or
								((vState = 498) and (hState = 476)) or
								((vState = 498) and (hState = 477)) or
								((vState = 498) and (hState = 478)) or
								((vState = 498) and (hState = 479)) or
								((vState = 498) and (hState = 480)) or
								((vState = 498) and (hState = 522)) or
								((vState = 498) and (hState = 536)) or
								((vState = 498) and (hState = 537)) or
								((vState = 498) and (hState = 538)) or
								((vState = 498) and (hState = 539)) or
								((vState = 498) and (hState = 540)) or
								((vState = 498) and (hState = 541)) or
								((vState = 498) and (hState = 542)) or
								((vState = 498) and (hState = 543)) or
								((vState = 498) and (hState = 544)) or
								((vState = 498) and (hState = 545)) or
								((vState = 498) and (hState = 546)) or
								((vState = 498) and (hState = 547)) or
								((vState = 498) and (hState = 548)) or
								((vState = 498) and (hState = 569)) or
								((vState = 498) and (hState = 570)) or
								((vState = 498) and (hState = 571)) or
								((vState = 498) and (hState = 572)) or
								((vState = 498) and (hState = 573)) or
								((vState = 498) and (hState = 574)) or
								((vState = 498) and (hState = 575)) or
								((vState = 498) and (hState = 576)) or
								((vState = 498) and (hState = 577)) or
								((vState = 498) and (hState = 578)) or
								((vState = 498) and (hState = 579)) or
								((vState = 498) and (hState = 580)) or
								((vState = 498) and (hState = 581)) or
								((vState = 498) and (hState = 582)) or
								((vState = 498) and (hState = 583)) or
								((vState = 498) and (hState = 584)) or
								((vState = 498) and (hState = 585)) or
								((vState = 498) and (hState = 586)) or
								((vState = 498) and (hState = 587)) or
								((vState = 498) and (hState = 588)) or
								((vState = 498) and (hState = 589)) or
								((vState = 498) and (hState = 590)) or
								((vState = 498) and (hState = 591)) or
								((vState = 498) and (hState = 592)) or
								((vState = 498) and (hState = 593)) or
								((vState = 498) and (hState = 594)) or
								((vState = 498) and (hState = 595)) or
								((vState = 498) and (hState = 596)) or
								((vState = 498) and (hState = 597)) or
								((vState = 499) and (hState = 319)) or
								((vState = 499) and (hState = 331)) or
								((vState = 499) and (hState = 347)) or
								((vState = 499) and (hState = 363)) or
								((vState = 499) and (hState = 373)) or
								((vState = 499) and (hState = 374)) or
								((vState = 499) and (hState = 375)) or
								((vState = 499) and (hState = 383)) or
								((vState = 499) and (hState = 389)) or
								((vState = 499) and (hState = 453)) or
								((vState = 499) and (hState = 485)) or
								((vState = 499) and (hState = 502)) or
								((vState = 499) and (hState = 519)) or
								((vState = 499) and (hState = 537)) or
								((vState = 499) and (hState = 541)) or
								((vState = 499) and (hState = 542)) or
								((vState = 499) and (hState = 543)) or
								((vState = 499) and (hState = 544)) or
								((vState = 499) and (hState = 545)) or
								((vState = 499) and (hState = 546)) or
								((vState = 499) and (hState = 547)) or
								((vState = 499) and (hState = 548)) or
								((vState = 499) and (hState = 549)) or
								((vState = 499) and (hState = 550)) or
								((vState = 499) and (hState = 551)) or
								((vState = 499) and (hState = 552)) or
								((vState = 499) and (hState = 553)) or
								((vState = 499) and (hState = 554)) or
								((vState = 499) and (hState = 555)) or
								((vState = 499) and (hState = 556)) or
								((vState = 499) and (hState = 557)) or
								((vState = 499) and (hState = 558)) or
								((vState = 499) and (hState = 559)) or
								((vState = 499) and (hState = 560)) or
								((vState = 499) and (hState = 561)) or
								((vState = 499) and (hState = 562)) or
								((vState = 499) and (hState = 563)) or
								((vState = 499) and (hState = 564)) or
								((vState = 499) and (hState = 565)) or
								((vState = 499) and (hState = 566)) or
								((vState = 499) and (hState = 567)) or
								((vState = 499) and (hState = 568)) or
								((vState = 499) and (hState = 569)) or
								((vState = 499) and (hState = 570)) or
								((vState = 499) and (hState = 574)) or
								((vState = 499) and (hState = 575)) or
								((vState = 499) and (hState = 576)) or
								((vState = 499) and (hState = 577)) or
								((vState = 499) and (hState = 583)) or
								((vState = 499) and (hState = 584)) or
								((vState = 499) and (hState = 590)) or
								((vState = 499) and (hState = 591)) or
								((vState = 499) and (hState = 592)) or
								((vState = 499) and (hState = 593)) or
								((vState = 499) and (hState = 594)) or
								((vState = 499) and (hState = 595)) or
								((vState = 500) and (hState = 320)) or
								((vState = 500) and (hState = 345)) or
								((vState = 500) and (hState = 373)) or
								((vState = 500) and (hState = 383)) or
								((vState = 500) and (hState = 386)) or
								((vState = 500) and (hState = 387)) or
								((vState = 500) and (hState = 455)) or
								((vState = 500) and (hState = 501)) or
								((vState = 500) and (hState = 518)) or
								((vState = 500) and (hState = 537)) or
								((vState = 500) and (hState = 546)) or
								((vState = 500) and (hState = 563)) or
								((vState = 500) and (hState = 564)) or
								((vState = 500) and (hState = 565)) or
								((vState = 500) and (hState = 566)) or
								((vState = 500) and (hState = 567)) or
								((vState = 500) and (hState = 568)) or
								((vState = 500) and (hState = 569)) or
								((vState = 500) and (hState = 570)) or
								((vState = 500) and (hState = 574)) or
								((vState = 500) and (hState = 575)) or
								((vState = 500) and (hState = 576)) or
								((vState = 500) and (hState = 577)) or
								((vState = 500) and (hState = 583)) or
								((vState = 500) and (hState = 584)) or
								((vState = 500) and (hState = 590)) or
								((vState = 500) and (hState = 591)) or
								((vState = 500) and (hState = 592)) or
								((vState = 500) and (hState = 593)) or
								((vState = 501) and (hState = 383)) or
								((vState = 501) and (hState = 567)) or
								((vState = 501) and (hState = 568)) or
								((vState = 501) and (hState = 569)) or
								((vState = 501) and (hState = 570)) or
								((vState = 501) and (hState = 574)) or
								((vState = 501) and (hState = 575)) or
								((vState = 501) and (hState = 576)) or
								((vState = 501) and (hState = 577)) or
								((vState = 501) and (hState = 583)) or
								((vState = 501) and (hState = 590)) or
								((vState = 501) and (hState = 591)) or
								((vState = 502) and (hState = 383)) or
								((vState = 502) and (hState = 384)) or
								((vState = 502) and (hState = 572)) or
								((vState = 502) and (hState = 582)) or
								((vState = 502) and (hState = 583)) or
								((vState = 502) and (hState = 589)) or
								((vState = 503) and (hState = 335)) or
								((vState = 503) and (hState = 340)) or
								((vState = 503) and (hState = 366)) or
								((vState = 503) and (hState = 367)) or
								((vState = 503) and (hState = 368)) or
								((vState = 503) and (hState = 383)) or
								((vState = 503) and (hState = 384)) or
								((vState = 503) and (hState = 459)) or
								((vState = 503) and (hState = 460)) or
								((vState = 503) and (hState = 487)) or
								((vState = 503) and (hState = 497)) or
								((vState = 503) and (hState = 513)) or
								((vState = 503) and (hState = 536)) or
								((vState = 503) and (hState = 572)) or
								((vState = 503) and (hState = 582)) or
								((vState = 503) and (hState = 583)) or
								((vState = 503) and (hState = 588)) or
								((vState = 503) and (hState = 589)) or
								((vState = 504) and (hState = 336)) or
								((vState = 504) and (hState = 337)) or
								((vState = 504) and (hState = 338)) or
								((vState = 504) and (hState = 366)) or
								((vState = 504) and (hState = 367)) or
								((vState = 504) and (hState = 382)) or
								((vState = 504) and (hState = 383)) or
								((vState = 504) and (hState = 512)) or
								((vState = 504) and (hState = 536)) or
								((vState = 504) and (hState = 572)) or
								((vState = 504) and (hState = 582)) or
								((vState = 504) and (hState = 583)) or
								((vState = 504) and (hState = 584)) or
								((vState = 504) and (hState = 585)) or
								((vState = 504) and (hState = 586)) or
								((vState = 504) and (hState = 587)) or
								((vState = 504) and (hState = 588)) or
								((vState = 505) and (hState = 324)) or
								((vState = 505) and (hState = 363)) or
								((vState = 505) and (hState = 364)) or
								((vState = 505) and (hState = 365)) or
								((vState = 505) and (hState = 366)) or
								((vState = 505) and (hState = 367)) or
								((vState = 505) and (hState = 395)) or
								((vState = 505) and (hState = 464)) or
								((vState = 505) and (hState = 490)) or
								((vState = 505) and (hState = 536)) or
								((vState = 505) and (hState = 582)) or
								((vState = 505) and (hState = 583)) or
								((vState = 505) and (hState = 584)) or
								((vState = 505) and (hState = 585)) or
								((vState = 505) and (hState = 586)) or
								((vState = 505) and (hState = 587)) or
								((vState = 505) and (hState = 588)) or
								((vState = 506) and (hState = 509)) or
								((vState = 506) and (hState = 582)) or
								((vState = 506) and (hState = 583)) or
								((vState = 506) and (hState = 584)) or
								((vState = 507) and (hState = 368)) or
								((vState = 507) and (hState = 384)) or
								((vState = 507) and (hState = 507)) or
								((vState = 507) and (hState = 508)) or
								((vState = 507) and (hState = 509)) or
								((vState = 507) and (hState = 582)) or
								((vState = 507) and (hState = 583)) or
								((vState = 508) and (hState = 336)) or
								((vState = 508) and (hState = 337)) or
								((vState = 508) and (hState = 338)) or
								((vState = 508) and (hState = 339)) or
								((vState = 508) and (hState = 340)) or
								((vState = 508) and (hState = 341)) or
								((vState = 508) and (hState = 342)) or
								((vState = 508) and (hState = 343)) or
								((vState = 508) and (hState = 358)) or
								((vState = 508) and (hState = 359)) or
								((vState = 508) and (hState = 368)) or
								((vState = 508) and (hState = 377)) or
								((vState = 508) and (hState = 384)) or
								((vState = 508) and (hState = 392)) or
								((vState = 508) and (hState = 469)) or
								((vState = 508) and (hState = 492)) or
								((vState = 508) and (hState = 507)) or
								((vState = 508) and (hState = 508)) or
								((vState = 508) and (hState = 509)) or
								((vState = 508) and (hState = 510)) or
								((vState = 508) and (hState = 511)) or
								((vState = 508) and (hState = 512)) or
								((vState = 508) and (hState = 535)) or
								((vState = 508) and (hState = 541)) or
								((vState = 508) and (hState = 581)) or
								((vState = 508) and (hState = 582)) or
								((vState = 508) and (hState = 583)) or
								((vState = 508) and (hState = 592)) or
								((vState = 508) and (hState = 593)) or
								((vState = 509) and (hState = 346)) or
								((vState = 509) and (hState = 347)) or
								((vState = 509) and (hState = 348)) or
								((vState = 509) and (hState = 349)) or
								((vState = 509) and (hState = 350)) or
								((vState = 509) and (hState = 351)) or
								((vState = 509) and (hState = 352)) or
								((vState = 509) and (hState = 353)) or
								((vState = 509) and (hState = 354)) or
								((vState = 509) and (hState = 355)) or
								((vState = 509) and (hState = 356)) or
								((vState = 509) and (hState = 357)) or
								((vState = 509) and (hState = 384)) or
								((vState = 509) and (hState = 391)) or
								((vState = 509) and (hState = 470)) or
								((vState = 509) and (hState = 471)) or
								((vState = 509) and (hState = 516)) or
								((vState = 509) and (hState = 517)) or
								((vState = 509) and (hState = 518)) or
								((vState = 509) and (hState = 519)) or
								((vState = 509) and (hState = 535)) or
								((vState = 509) and (hState = 569)) or
								((vState = 509) and (hState = 579)) or
								((vState = 509) and (hState = 580)) or
								((vState = 509) and (hState = 581)) or
								((vState = 509) and (hState = 594)) or
								((vState = 509) and (hState = 595)) or
								((vState = 510) and (hState = 384)) or
								((vState = 510) and (hState = 390)) or
								((vState = 510) and (hState = 473)) or
								((vState = 510) and (hState = 474)) or
								((vState = 510) and (hState = 501)) or
								((vState = 510) and (hState = 523)) or
								((vState = 510) and (hState = 524)) or
								((vState = 510) and (hState = 525)) or
								((vState = 510) and (hState = 526)) or
								((vState = 510) and (hState = 527)) or
								((vState = 510) and (hState = 540)) or
								((vState = 510) and (hState = 577)) or
								((vState = 510) and (hState = 578)) or
								((vState = 510) and (hState = 579)) or
								((vState = 510) and (hState = 580)) or
								((vState = 510) and (hState = 581)) or
								((vState = 510) and (hState = 597)) or
								((vState = 511) and (hState = 384)) or
								((vState = 511) and (hState = 523)) or
								((vState = 511) and (hState = 524)) or
								((vState = 511) and (hState = 525)) or
								((vState = 511) and (hState = 526)) or
								((vState = 511) and (hState = 527)) or
								((vState = 511) and (hState = 540)) or
								((vState = 511) and (hState = 577)) or
								((vState = 511) and (hState = 578)) or
								((vState = 511) and (hState = 579)) or
								((vState = 511) and (hState = 580)) or
								((vState = 511) and (hState = 597)) or
								((vState = 511) and (hState = 598)) or
								((vState = 512) and (hState = 384)) or
								((vState = 512) and (hState = 523)) or
								((vState = 512) and (hState = 524)) or
								((vState = 512) and (hState = 525)) or
								((vState = 512) and (hState = 526)) or
								((vState = 512) and (hState = 527)) or
								((vState = 512) and (hState = 528)) or
								((vState = 512) and (hState = 529)) or
								((vState = 512) and (hState = 530)) or
								((vState = 512) and (hState = 531)) or
								((vState = 512) and (hState = 532)) or
								((vState = 512) and (hState = 533)) or
								((vState = 512) and (hState = 534)) or
								((vState = 512) and (hState = 539)) or
								((vState = 512) and (hState = 540)) or
								((vState = 512) and (hState = 577)) or
								((vState = 512) and (hState = 578)) or
								((vState = 512) and (hState = 579)) or
								((vState = 512) and (hState = 580)) or
								((vState = 512) and (hState = 597)) or
								((vState = 512) and (hState = 598)) or
								((vState = 512) and (hState = 599)) or
								((vState = 513) and (hState = 384)) or
								((vState = 513) and (hState = 528)) or
								((vState = 513) and (hState = 529)) or
								((vState = 513) and (hState = 530)) or
								((vState = 513) and (hState = 531)) or
								((vState = 513) and (hState = 532)) or
								((vState = 513) and (hState = 533)) or
								((vState = 513) and (hState = 534)) or
								((vState = 513) and (hState = 535)) or
								((vState = 513) and (hState = 536)) or
								((vState = 513) and (hState = 537)) or
								((vState = 513) and (hState = 538)) or
								((vState = 513) and (hState = 539)) or
								((vState = 513) and (hState = 540)) or
								((vState = 513) and (hState = 541)) or
								((vState = 513) and (hState = 577)) or
								((vState = 513) and (hState = 578)) or
								((vState = 513) and (hState = 579)) or
								((vState = 513) and (hState = 580)) or
								((vState = 514) and (hState = 384)) or
								((vState = 514) and (hState = 385)) or
								((vState = 514) and (hState = 386)) or
								((vState = 514) and (hState = 387)) or
								((vState = 514) and (hState = 480)) or
								((vState = 514) and (hState = 497)) or
								((vState = 514) and (hState = 506)) or
								((vState = 514) and (hState = 529)) or
								((vState = 514) and (hState = 530)) or
								((vState = 514) and (hState = 531)) or
								((vState = 514) and (hState = 532)) or
								((vState = 514) and (hState = 533)) or
								((vState = 514) and (hState = 534)) or
								((vState = 514) and (hState = 535)) or
								((vState = 514) and (hState = 536)) or
								((vState = 514) and (hState = 537)) or
								((vState = 514) and (hState = 538)) or
								((vState = 514) and (hState = 539)) or
								((vState = 514) and (hState = 540)) or
								((vState = 514) and (hState = 541)) or
								((vState = 514) and (hState = 542)) or
								((vState = 514) and (hState = 543)) or
								((vState = 514) and (hState = 544)) or
								((vState = 514) and (hState = 545)) or
								((vState = 514) and (hState = 546)) or
								((vState = 514) and (hState = 547)) or
								((vState = 514) and (hState = 548)) or
								((vState = 514) and (hState = 567)) or
								((vState = 514) and (hState = 577)) or
								((vState = 514) and (hState = 578)) or
								((vState = 514) and (hState = 579)) or
								((vState = 514) and (hState = 580)) or
								((vState = 514) and (hState = 588)) or
								((vState = 514) and (hState = 589)) or
								((vState = 514) and (hState = 590)) or
								((vState = 514) and (hState = 591)) or
								((vState = 515) and (hState = 384)) or
								((vState = 515) and (hState = 385)) or
								((vState = 515) and (hState = 482)) or
								((vState = 515) and (hState = 507)) or
								((vState = 515) and (hState = 532)) or
								((vState = 515) and (hState = 566)) or
								((vState = 515) and (hState = 567)) or
								((vState = 515) and (hState = 568)) or
								((vState = 515) and (hState = 569)) or
								((vState = 515) and (hState = 576)) or
								((vState = 515) and (hState = 577)) or
								((vState = 515) and (hState = 578)) or
								((vState = 515) and (hState = 579)) or
								((vState = 515) and (hState = 580)) or
								((vState = 515) and (hState = 581)) or
								((vState = 515) and (hState = 582)) or
								((vState = 515) and (hState = 583)) or
								((vState = 515) and (hState = 584)) or
								((vState = 516) and (hState = 532)) or
								((vState = 516) and (hState = 566)) or
								((vState = 516) and (hState = 567)) or
								((vState = 516) and (hState = 568)) or
								((vState = 516) and (hState = 569)) or
								((vState = 516) and (hState = 575)) or
								((vState = 516) and (hState = 576)) or
								((vState = 516) and (hState = 577)) or
								((vState = 516) and (hState = 578)) or
								((vState = 516) and (hState = 579)) or
								((vState = 517) and (hState = 532)) or
								((vState = 517) and (hState = 566)) or
								((vState = 517) and (hState = 567)) or
								((vState = 517) and (hState = 568)) or
								((vState = 517) and (hState = 569)) or
								((vState = 517) and (hState = 573)) or
								((vState = 517) and (hState = 579)) or
								((vState = 518) and (hState = 511)) or
								((vState = 518) and (hState = 532)) or
								((vState = 518) and (hState = 565)) or
								((vState = 518) and (hState = 571)) or
								((vState = 518) and (hState = 572)) or
								((vState = 518) and (hState = 579)) or
								((vState = 519) and (hState = 501)) or
								((vState = 519) and (hState = 512)) or
								((vState = 519) and (hState = 563)) or
								((vState = 519) and (hState = 564)) or
								((vState = 519) and (hState = 571)) or
								((vState = 519) and (hState = 572)) or
								((vState = 519) and (hState = 579)) or
								((vState = 520) and (hState = 502)) or
								((vState = 520) and (hState = 513)) or
								((vState = 520) and (hState = 531)) or
								((vState = 520) and (hState = 563)) or
								((vState = 520) and (hState = 579)) or
								((vState = 521) and (hState = 503)) or
								((vState = 521) and (hState = 514)) or
								((vState = 521) and (hState = 531)) or
								((vState = 521) and (hState = 563)) or
								((vState = 521) and (hState = 569)) or
								((vState = 521) and (hState = 579)) or
								((vState = 522) and (hState = 503)) or
								((vState = 522) and (hState = 531)) or
								((vState = 523) and (hState = 503)) or
								((vState = 524) and (hState = 490)) or
								((vState = 524) and (hState = 503)) or
								((vState = 524) and (hState = 518)) or
								((vState = 525) and (hState = 490)) or
								((vState = 525) and (hState = 519)) or
								((vState = 525) and (hState = 530)) or
								((vState = 526) and (hState = 530)) or
								((vState = 527) and (hState = 530)) or
								((vState = 528) and (hState = 491)) or
								((vState = 528) and (hState = 530)) or
								((vState = 529) and (hState = 491)) or
								((vState = 529) and (hState = 524)) or
								((vState = 529) and (hState = 530)) or
								((vState = 529) and (hState = 563)) or
								((vState = 529) and (hState = 583)) or
								((vState = 529) and (hState = 584)) or
								((vState = 529) and (hState = 585)) or
								((vState = 529) and (hState = 586)) or
								((vState = 529) and (hState = 587)) or
								((vState = 529) and (hState = 588)) or
								((vState = 530) and (hState = 525)) or
								((vState = 530) and (hState = 531)) or
								((vState = 530) and (hState = 558)) or
								((vState = 530) and (hState = 562)) or
								((vState = 530) and (hState = 574)) or
								((vState = 530) and (hState = 575)) or
								((vState = 530) and (hState = 576)) or
								((vState = 530) and (hState = 577)) or
								((vState = 530) and (hState = 578)) or
								((vState = 530) and (hState = 579)) or
								((vState = 531) and (hState = 492)) or
								((vState = 531) and (hState = 506)) or
								((vState = 531) and (hState = 532)) or
								((vState = 531) and (hState = 558)) or
								((vState = 531) and (hState = 559)) or
								((vState = 531) and (hState = 560)) or
								((vState = 531) and (hState = 561)) or
								((vState = 531) and (hState = 562)) or
								((vState = 531) and (hState = 567)) or
								((vState = 531) and (hState = 568)) or
								((vState = 531) and (hState = 569)) or
								((vState = 531) and (hState = 570)) or
								((vState = 531) and (hState = 571)) or
								((vState = 531) and (hState = 572)) or
								((vState = 532) and (hState = 492)) or
								((vState = 532) and (hState = 506)) or
								((vState = 532) and (hState = 558)) or
								((vState = 532) and (hState = 559)) or
								((vState = 532) and (hState = 560)) or
								((vState = 532) and (hState = 561)) or
								((vState = 532) and (hState = 562)) or
								((vState = 533) and (hState = 492)) or
								((vState = 533) and (hState = 506)) or
								((vState = 533) and (hState = 557)) or
								((vState = 533) and (hState = 558)) or
								((vState = 533) and (hState = 595)) or
								((vState = 534) and (hState = 506)) or
								((vState = 534) and (hState = 535)) or
								((vState = 534) and (hState = 554)) or
								((vState = 534) and (hState = 555)) or
								((vState = 534) and (hState = 556)) or
								((vState = 534) and (hState = 557)) or
								((vState = 535) and (hState = 531)) or
								((vState = 535) and (hState = 535)) or
								((vState = 535) and (hState = 536)) or
								((vState = 535) and (hState = 542)) or
								((vState = 535) and (hState = 543)) or
								((vState = 535) and (hState = 544)) or
								((vState = 535) and (hState = 545)) or
								((vState = 535) and (hState = 546)) or
								((vState = 535) and (hState = 547)) or
								((vState = 535) and (hState = 548)) or
								((vState = 535) and (hState = 555)) or
								((vState = 535) and (hState = 556)) or
								((vState = 535) and (hState = 557)) or
								((vState = 536) and (hState = 507)) or
								((vState = 536) and (hState = 534)) or
								((vState = 536) and (hState = 535)) or
								((vState = 536) and (hState = 536)) or
								((vState = 536) and (hState = 537)) or
								((vState = 536) and (hState = 542)) or
								((vState = 536) and (hState = 555)) or
								((vState = 536) and (hState = 556)) or
								((vState = 536) and (hState = 594)) or
								((vState = 537) and (hState = 507)) or
								((vState = 537) and (hState = 535)) or
								((vState = 537) and (hState = 536)) or
								((vState = 537) and (hState = 537)) or
								((vState = 537) and (hState = 538)) or
								((vState = 537) and (hState = 594)) or
								((vState = 538) and (hState = 507)) or
								((vState = 538) and (hState = 536)) or
								((vState = 538) and (hState = 537)) or
								((vState = 538) and (hState = 538)) or
								((vState = 538) and (hState = 539)) or
								((vState = 539) and (hState = 537)) or
								((vState = 539) and (hState = 538)) or
								((vState = 539) and (hState = 539)) or
								((vState = 539) and (hState = 540)) or
								((vState = 539) and (hState = 544)) or
								((vState = 539) and (hState = 568)) or
								((vState = 540) and (hState = 537)) or
								((vState = 540) and (hState = 538)) or
								((vState = 540) and (hState = 539)) or
								((vState = 540) and (hState = 540)) or
								((vState = 540) and (hState = 541)) or
								((vState = 540) and (hState = 542)) or
								((vState = 540) and (hState = 543)) or
								((vState = 540) and (hState = 544)) or
								((vState = 540) and (hState = 566)) or
								((vState = 540) and (hState = 567)) or
								((vState = 540) and (hState = 568)) or
								((vState = 540) and (hState = 593)) or
								((vState = 541) and (hState = 508)) or
								((vState = 541) and (hState = 540)) or
								((vState = 541) and (hState = 541)) or
								((vState = 541) and (hState = 542)) or
								((vState = 541) and (hState = 543)) or
								((vState = 541) and (hState = 544)) or
								((vState = 541) and (hState = 545)) or
								((vState = 541) and (hState = 563)) or
								((vState = 541) and (hState = 564)) or
								((vState = 541) and (hState = 565)) or
								((vState = 541) and (hState = 593)) or
								((vState = 542) and (hState = 508)) or
								((vState = 542) and (hState = 541)) or
								((vState = 542) and (hState = 542)) or
								((vState = 542) and (hState = 543)) or
								((vState = 542) and (hState = 544)) or
								((vState = 542) and (hState = 545)) or
								((vState = 542) and (hState = 546)) or
								((vState = 542) and (hState = 562)) or
								((vState = 542) and (hState = 563)) or
								((vState = 542) and (hState = 564)) or
								((vState = 542) and (hState = 583)) or
								((vState = 543) and (hState = 508)) or
								((vState = 543) and (hState = 542)) or
								((vState = 543) and (hState = 543)) or
								((vState = 543) and (hState = 544)) or
								((vState = 543) and (hState = 545)) or
								((vState = 543) and (hState = 546)) or
								((vState = 543) and (hState = 562)) or
								((vState = 543) and (hState = 563)) or
								((vState = 544) and (hState = 496)) or
								((vState = 544) and (hState = 544)) or
								((vState = 544) and (hState = 545)) or
								((vState = 544) and (hState = 546)) or
								((vState = 544) and (hState = 547)) or
								((vState = 544) and (hState = 560)) or
								((vState = 544) and (hState = 561)) or
								((vState = 544) and (hState = 580)) or
								((vState = 544) and (hState = 581)) or
								((vState = 545) and (hState = 496)) or
								((vState = 545) and (hState = 529)) or
								((vState = 545) and (hState = 530)) or
								((vState = 545) and (hState = 544)) or
								((vState = 545) and (hState = 545)) or
								((vState = 545) and (hState = 546)) or
								((vState = 545) and (hState = 547)) or
								((vState = 545) and (hState = 557)) or
								((vState = 545) and (hState = 558)) or
								((vState = 545) and (hState = 559)) or
								((vState = 545) and (hState = 560)) or
								((vState = 545) and (hState = 579)) or
								((vState = 545) and (hState = 580)) or
								((vState = 545) and (hState = 581)) or
								((vState = 546) and (hState = 529)) or
								((vState = 546) and (hState = 530)) or
								((vState = 546) and (hState = 546)) or
								((vState = 546) and (hState = 547)) or
								((vState = 546) and (hState = 548)) or
								((vState = 546) and (hState = 558)) or
								((vState = 546) and (hState = 559)) or
								((vState = 546) and (hState = 577)) or
								((vState = 546) and (hState = 578)) or
								((vState = 546) and (hState = 579)) or
								((vState = 546) and (hState = 580)) or
								((vState = 546) and (hState = 597)) or
								((vState = 547) and (hState = 497)) or
								((vState = 547) and (hState = 528)) or
								((vState = 547) and (hState = 529)) or
								((vState = 547) and (hState = 530)) or
								((vState = 547) and (hState = 547)) or
								((vState = 547) and (hState = 548)) or
								((vState = 547) and (hState = 549)) or
								((vState = 547) and (hState = 550)) or
								((vState = 547) and (hState = 551)) or
								((vState = 547) and (hState = 552)) or
								((vState = 547) and (hState = 558)) or
								((vState = 547) and (hState = 579)) or
								((vState = 547) and (hState = 580)) or
								((vState = 547) and (hState = 590)) or
								((vState = 547) and (hState = 594)) or
								((vState = 547) and (hState = 595)) or
								((vState = 547) and (hState = 596)) or
								((vState = 548) and (hState = 497)) or
								((vState = 548) and (hState = 527)) or
								((vState = 548) and (hState = 530)) or
								((vState = 548) and (hState = 547)) or
								((vState = 548) and (hState = 548)) or
								((vState = 548) and (hState = 549)) or
								((vState = 548) and (hState = 550)) or
								((vState = 548) and (hState = 551)) or
								((vState = 548) and (hState = 579)) or
								((vState = 548) and (hState = 590)) or
								((vState = 548) and (hState = 594)) or
								((vState = 548) and (hState = 595)) or
								((vState = 549) and (hState = 497)) or
								((vState = 549) and (hState = 527)) or
								((vState = 549) and (hState = 530)) or
								((vState = 549) and (hState = 547)) or
								((vState = 549) and (hState = 548)) or
								((vState = 549) and (hState = 549)) or
								((vState = 549) and (hState = 550)) or
								((vState = 549) and (hState = 551)) or
								((vState = 549) and (hState = 590)) or
								((vState = 549) and (hState = 591)) or
								((vState = 549) and (hState = 592)) or
								((vState = 549) and (hState = 593)) or
								((vState = 549) and (hState = 594)) or
								((vState = 550) and (hState = 497)) or
								((vState = 550) and (hState = 526)) or
								((vState = 550) and (hState = 527)) or
								((vState = 550) and (hState = 530)) or
								((vState = 550) and (hState = 547)) or
								((vState = 550) and (hState = 548)) or
								((vState = 550) and (hState = 549)) or
								((vState = 550) and (hState = 550)) or
								((vState = 550) and (hState = 551)) or
								((vState = 550) and (hState = 571)) or
								((vState = 550) and (hState = 572)) or
								((vState = 550) and (hState = 590)) or
								((vState = 550) and (hState = 591)) or
								((vState = 550) and (hState = 592)) or
								((vState = 550) and (hState = 593)) or
								((vState = 550) and (hState = 594)) or
								((vState = 551) and (hState = 511)) or
								((vState = 551) and (hState = 525)) or
								((vState = 551) and (hState = 551)) or
								((vState = 551) and (hState = 552)) or
								((vState = 551) and (hState = 553)) or
								((vState = 551) and (hState = 569)) or
								((vState = 551) and (hState = 570)) or
								((vState = 551) and (hState = 571)) or
								((vState = 551) and (hState = 572)) or
								((vState = 551) and (hState = 578)) or
								((vState = 551) and (hState = 590)) or
								((vState = 551) and (hState = 591)) or
								((vState = 551) and (hState = 592)) or
								((vState = 551) and (hState = 593)) or
								((vState = 551) and (hState = 594)) or
								((vState = 552) and (hState = 511)) or
								((vState = 552) and (hState = 542)) or
								((vState = 552) and (hState = 551)) or
								((vState = 552) and (hState = 552)) or
								((vState = 552) and (hState = 553)) or
								((vState = 552) and (hState = 568)) or
								((vState = 552) and (hState = 569)) or
								((vState = 552) and (hState = 570)) or
								((vState = 552) and (hState = 571)) or
								((vState = 552) and (hState = 572)) or
								((vState = 552) and (hState = 577)) or
								((vState = 552) and (hState = 589)) or
								((vState = 552) and (hState = 593)) or
								((vState = 553) and (hState = 511)) or
								((vState = 553) and (hState = 553)) or
								((vState = 553) and (hState = 554)) or
								((vState = 553) and (hState = 568)) or
								((vState = 553) and (hState = 577)) or
								((vState = 553) and (hState = 589)) or
								((vState = 554) and (hState = 531)) or
								((vState = 554) and (hState = 555)) or
								((vState = 554) and (hState = 567)) or
								((vState = 554) and (hState = 568)) or
								((vState = 554) and (hState = 588)) or
								((vState = 554) and (hState = 589)) or
								((vState = 555) and (hState = 531)) or
								((vState = 555) and (hState = 537)) or
								((vState = 555) and (hState = 548)) or
								((vState = 555) and (hState = 555)) or
								((vState = 555) and (hState = 556)) or
								((vState = 555) and (hState = 557)) or
								((vState = 555) and (hState = 564)) or
								((vState = 555) and (hState = 565)) or
								((vState = 555) and (hState = 566)) or
								((vState = 555) and (hState = 567)) or
								((vState = 555) and (hState = 568)) or
								((vState = 555) and (hState = 574)) or
								((vState = 555) and (hState = 575)) or
								((vState = 555) and (hState = 588)) or
								((vState = 555) and (hState = 589)) or
								((vState = 555) and (hState = 590)) or
								((vState = 556) and (hState = 512)) or
								((vState = 556) and (hState = 531)) or
								((vState = 556) and (hState = 535)) or
								((vState = 556) and (hState = 536)) or
								((vState = 556) and (hState = 537)) or
								((vState = 556) and (hState = 538)) or
								((vState = 556) and (hState = 547)) or
								((vState = 556) and (hState = 555)) or
								((vState = 556) and (hState = 556)) or
								((vState = 556) and (hState = 557)) or
								((vState = 556) and (hState = 558)) or
								((vState = 556) and (hState = 559)) or
								((vState = 556) and (hState = 563)) or
								((vState = 556) and (hState = 564)) or
								((vState = 556) and (hState = 565)) or
								((vState = 556) and (hState = 566)) or
								((vState = 556) and (hState = 567)) or
								((vState = 556) and (hState = 568)) or
								((vState = 556) and (hState = 574)) or
								((vState = 556) and (hState = 575)) or
								((vState = 556) and (hState = 584)) or
								((vState = 556) and (hState = 588)) or
								((vState = 556) and (hState = 589)) or
								((vState = 556) and (hState = 590)) or
								((vState = 557) and (hState = 512)) or
								((vState = 557) and (hState = 522)) or
								((vState = 557) and (hState = 525)) or
								((vState = 557) and (hState = 526)) or
								((vState = 557) and (hState = 527)) or
								((vState = 557) and (hState = 528)) or
								((vState = 557) and (hState = 529)) or
								((vState = 557) and (hState = 530)) or
								((vState = 557) and (hState = 531)) or
								((vState = 557) and (hState = 532)) or
								((vState = 557) and (hState = 533)) or
								((vState = 557) and (hState = 534)) or
								((vState = 557) and (hState = 535)) or
								((vState = 557) and (hState = 536)) or
								((vState = 557) and (hState = 537)) or
								((vState = 557) and (hState = 538)) or
								((vState = 557) and (hState = 539)) or
								((vState = 557) and (hState = 540)) or
								((vState = 557) and (hState = 541)) or
								((vState = 557) and (hState = 542)) or
								((vState = 557) and (hState = 543)) or
								((vState = 557) and (hState = 544)) or
								((vState = 557) and (hState = 545)) or
								((vState = 557) and (hState = 546)) or
								((vState = 557) and (hState = 547)) or
								((vState = 557) and (hState = 555)) or
								((vState = 557) and (hState = 556)) or
								((vState = 557) and (hState = 557)) or
								((vState = 557) and (hState = 558)) or
								((vState = 557) and (hState = 559)) or
								((vState = 557) and (hState = 560)) or
								((vState = 557) and (hState = 561)) or
								((vState = 557) and (hState = 562)) or
								((vState = 557) and (hState = 563)) or
								((vState = 557) and (hState = 564)) or
								((vState = 557) and (hState = 565)) or
								((vState = 557) and (hState = 566)) or
								((vState = 557) and (hState = 567)) or
								((vState = 557) and (hState = 568)) or
								((vState = 557) and (hState = 569)) or
								((vState = 557) and (hState = 570)) or
								((vState = 557) and (hState = 571)) or
								((vState = 557) and (hState = 572)) or
								((vState = 557) and (hState = 573)) or
								((vState = 557) and (hState = 574)) or
								((vState = 557) and (hState = 575)) or
								((vState = 557) and (hState = 576)) or
								((vState = 557) and (hState = 577)) or
								((vState = 557) and (hState = 578)) or
								((vState = 557) and (hState = 579)) or
								((vState = 557) and (hState = 580)) or
								((vState = 557) and (hState = 581)) or
								((vState = 557) and (hState = 582)) or
								((vState = 557) and (hState = 583)) or
								((vState = 557) and (hState = 584)) or
								((vState = 557) and (hState = 588)) or
								((vState = 557) and (hState = 589)) or
								((vState = 558) and (hState = 511)) or
								((vState = 558) and (hState = 512)) or
								((vState = 558) and (hState = 513)) or
								((vState = 558) and (hState = 521)) or
								((vState = 558) and (hState = 522)) or
								((vState = 558) and (hState = 530)) or
								((vState = 558) and (hState = 531)) or
								((vState = 558) and (hState = 532)) or
								((vState = 558) and (hState = 533)) or
								((vState = 558) and (hState = 534)) or
								((vState = 558) and (hState = 535)) or
								((vState = 558) and (hState = 536)) or
								((vState = 558) and (hState = 537)) or
								((vState = 558) and (hState = 538)) or
								((vState = 558) and (hState = 539)) or
								((vState = 558) and (hState = 540)) or
								((vState = 558) and (hState = 541)) or
								((vState = 558) and (hState = 542)) or
								((vState = 558) and (hState = 543)) or
								((vState = 558) and (hState = 544)) or
								((vState = 558) and (hState = 545)) or
								((vState = 558) and (hState = 546)) or
								((vState = 558) and (hState = 547)) or
								((vState = 558) and (hState = 548)) or
								((vState = 558) and (hState = 554)) or
								((vState = 558) and (hState = 555)) or
								((vState = 558) and (hState = 556)) or
								((vState = 558) and (hState = 557)) or
								((vState = 558) and (hState = 558)) or
								((vState = 558) and (hState = 559)) or
								((vState = 558) and (hState = 563)) or
								((vState = 558) and (hState = 564)) or
								((vState = 558) and (hState = 565)) or
								((vState = 558) and (hState = 573)) or
								((vState = 558) and (hState = 578)) or
								((vState = 558) and (hState = 579)) or
								((vState = 558) and (hState = 580)) or
								((vState = 558) and (hState = 581)) or
								((vState = 558) and (hState = 588)) or
								((vState = 559) and (hState = 499)) or
								((vState = 559) and (hState = 500)) or
								((vState = 559) and (hState = 513)) or
								((vState = 559) and (hState = 519)) or
								((vState = 559) and (hState = 520)) or
								((vState = 559) and (hState = 532)) or
								((vState = 559) and (hState = 533)) or
								((vState = 559) and (hState = 540)) or
								((vState = 559) and (hState = 541)) or
								((vState = 559) and (hState = 542)) or
								((vState = 559) and (hState = 546)) or
								((vState = 559) and (hState = 547)) or
								((vState = 559) and (hState = 556)) or
								((vState = 559) and (hState = 557)) or
								((vState = 559) and (hState = 558)) or
								((vState = 559) and (hState = 559)) or
								((vState = 559) and (hState = 578)) or
								((vState = 559) and (hState = 579)) or
								((vState = 559) and (hState = 580)) or
								((vState = 559) and (hState = 588)) or
								((vState = 560) and (hState = 487)) or
								((vState = 560) and (hState = 488)) or
								((vState = 560) and (hState = 501)) or
								((vState = 560) and (hState = 513)) or
								((vState = 560) and (hState = 519)) or
								((vState = 560) and (hState = 532)) or
								((vState = 560) and (hState = 540)) or
								((vState = 560) and (hState = 547)) or
								((vState = 560) and (hState = 556)) or
								((vState = 560) and (hState = 557)) or
								((vState = 560) and (hState = 558)) or
								((vState = 560) and (hState = 559)) or
								((vState = 560) and (hState = 560)) or
								((vState = 560) and (hState = 578)) or
								((vState = 560) and (hState = 579)) or
								((vState = 560) and (hState = 580)) or
								((vState = 560) and (hState = 587)) or
								((vState = 561) and (hState = 487)) or
								((vState = 561) and (hState = 488)) or
								((vState = 561) and (hState = 501)) or
								((vState = 561) and (hState = 513)) or
								((vState = 561) and (hState = 519)) or
								((vState = 561) and (hState = 532)) or
								((vState = 561) and (hState = 540)) or
								((vState = 561) and (hState = 547)) or
								((vState = 561) and (hState = 556)) or
								((vState = 561) and (hState = 557)) or
								((vState = 561) and (hState = 558)) or
								((vState = 561) and (hState = 559)) or
								((vState = 561) and (hState = 560)) or
								((vState = 561) and (hState = 561)) or
								((vState = 561) and (hState = 568)) or
								((vState = 561) and (hState = 572)) or
								((vState = 561) and (hState = 576)) or
								((vState = 561) and (hState = 577)) or
								((vState = 561) and (hState = 578)) or
								((vState = 561) and (hState = 579)) or
								((vState = 561) and (hState = 580)) or
								((vState = 561) and (hState = 595)) or
								((vState = 562) and (hState = 501)) or
								((vState = 562) and (hState = 513)) or
								((vState = 562) and (hState = 532)) or
								((vState = 562) and (hState = 548)) or
								((vState = 562) and (hState = 560)) or
								((vState = 562) and (hState = 561)) or
								((vState = 562) and (hState = 562)) or
								((vState = 562) and (hState = 563)) or
								((vState = 562) and (hState = 564)) or
								((vState = 562) and (hState = 569)) or
								((vState = 562) and (hState = 570)) or
								((vState = 562) and (hState = 571)) or
								((vState = 562) and (hState = 572)) or
								((vState = 562) and (hState = 573)) or
								((vState = 562) and (hState = 574)) or
								((vState = 562) and (hState = 575)) or
								((vState = 562) and (hState = 576)) or
								((vState = 562) and (hState = 577)) or
								((vState = 562) and (hState = 594)) or
								((vState = 562) and (hState = 595)) or
								((vState = 563) and (hState = 490)) or
								((vState = 563) and (hState = 502)) or
								((vState = 563) and (hState = 513)) or
								((vState = 563) and (hState = 518)) or
								((vState = 563) and (hState = 532)) or
								((vState = 563) and (hState = 537)) or
								((vState = 563) and (hState = 550)) or
								((vState = 563) and (hState = 551)) or
								((vState = 563) and (hState = 552)) or
								((vState = 563) and (hState = 560)) or
								((vState = 563) and (hState = 561)) or
								((vState = 563) and (hState = 562)) or
								((vState = 563) and (hState = 563)) or
								((vState = 563) and (hState = 564)) or
								((vState = 563) and (hState = 569)) or
								((vState = 563) and (hState = 570)) or
								((vState = 563) and (hState = 571)) or
								((vState = 563) and (hState = 572)) or
								((vState = 563) and (hState = 573)) or
								((vState = 563) and (hState = 574)) or
								((vState = 563) and (hState = 575)) or
								((vState = 563) and (hState = 584)) or
								((vState = 563) and (hState = 585)) or
								((vState = 563) and (hState = 594)) or
								((vState = 564) and (hState = 518)) or
								((vState = 564) and (hState = 532)) or
								((vState = 564) and (hState = 533)) or
								((vState = 564) and (hState = 550)) or
								((vState = 564) and (hState = 551)) or
								((vState = 564) and (hState = 552)) or
								((vState = 564) and (hState = 561)) or
								((vState = 564) and (hState = 562)) or
								((vState = 564) and (hState = 563)) or
								((vState = 564) and (hState = 564)) or
								((vState = 564) and (hState = 573)) or
								((vState = 564) and (hState = 574)) or
								((vState = 564) and (hState = 575)) or
								((vState = 564) and (hState = 584)) or
								((vState = 564) and (hState = 585)) or
								((vState = 565) and (hState = 532)) or
								((vState = 565) and (hState = 533)) or
								((vState = 565) and (hState = 534)) or
								((vState = 565) and (hState = 550)) or
								((vState = 565) and (hState = 562)) or
								((vState = 565) and (hState = 573)) or
								((vState = 565) and (hState = 574)) or
								((vState = 565) and (hState = 575)) or
								((vState = 565) and (hState = 576)) or
								((vState = 565) and (hState = 584)) or
								((vState = 565) and (hState = 585)) or
								((vState = 565) and (hState = 593)) or
								((vState = 566) and (hState = 492)) or
								((vState = 566) and (hState = 519)) or
								((vState = 566) and (hState = 532)) or
								((vState = 566) and (hState = 533)) or
								((vState = 566) and (hState = 553)) or
								((vState = 566) and (hState = 562)) or
								((vState = 566) and (hState = 566)) or
								((vState = 566) and (hState = 573)) or
								((vState = 566) and (hState = 574)) or
								((vState = 566) and (hState = 575)) or
								((vState = 566) and (hState = 576)) or
								((vState = 566) and (hState = 577)) or
								((vState = 566) and (hState = 583)) or
								((vState = 566) and (hState = 584)) or
								((vState = 566) and (hState = 585)) or
								((vState = 566) and (hState = 592)) or
								((vState = 566) and (hState = 593)) or
								((vState = 567) and (hState = 532)) or
								((vState = 567) and (hState = 533)) or
								((vState = 567) and (hState = 547)) or
								((vState = 567) and (hState = 562)) or
								((vState = 567) and (hState = 567)) or
								((vState = 567) and (hState = 572)) or
								((vState = 567) and (hState = 578)) or
								((vState = 567) and (hState = 583)) or
								((vState = 567) and (hState = 584)) or
								((vState = 567) and (hState = 588)) or
								((vState = 568) and (hState = 506)) or
								((vState = 568) and (hState = 522)) or
								((vState = 568) and (hState = 531)) or
								((vState = 568) and (hState = 532)) or
								((vState = 568) and (hState = 533)) or
								((vState = 568) and (hState = 546)) or
								((vState = 568) and (hState = 556)) or
								((vState = 568) and (hState = 562)) or
								((vState = 568) and (hState = 563)) or
								((vState = 568) and (hState = 568)) or
								((vState = 568) and (hState = 569)) or
								((vState = 568) and (hState = 570)) or
								((vState = 568) and (hState = 581)) or
								((vState = 568) and (hState = 582)) or
								((vState = 568) and (hState = 583)) or
								((vState = 568) and (hState = 584)) or
								((vState = 568) and (hState = 589)) or
								((vState = 568) and (hState = 590)) or
								((vState = 568) and (hState = 591)) or
								((vState = 569) and (hState = 568)) or
								((vState = 569) and (hState = 569)) or
								((vState = 569) and (hState = 570)) or
								((vState = 569) and (hState = 581)) or
								((vState = 569) and (hState = 582)) or
								((vState = 569) and (hState = 583)) or
								((vState = 569) and (hState = 584)) or
								((vState = 569) and (hState = 589)) or
								((vState = 569) and (hState = 590)) or
								((vState = 569) and (hState = 591)) or
								((vState = 570) and (hState = 560)) or
								((vState = 570) and (hState = 589)) or
								((vState = 570) and (hState = 590)) or
								((vState = 570) and (hState = 591)) or
								((vState = 571) and (hState = 496)) or
								((vState = 571) and (hState = 508)) or
								((vState = 571) and (hState = 524)) or
								((vState = 571) and (hState = 527)) or
								((vState = 571) and (hState = 528)) or
								((vState = 571) and (hState = 542)) or
								((vState = 571) and (hState = 560)) or
								((vState = 571) and (hState = 565)) or
								((vState = 571) and (hState = 566)) or
								((vState = 571) and (hState = 567)) or
								((vState = 571) and (hState = 571)) or
								((vState = 571) and (hState = 589)) or
								((vState = 571) and (hState = 590)) or
								((vState = 571) and (hState = 591)) or
								((vState = 572) and (hState = 497)) or
								((vState = 572) and (hState = 524)) or
								((vState = 572) and (hState = 525)) or
								((vState = 572) and (hState = 526)) or
								((vState = 572) and (hState = 527)) or
								((vState = 572) and (hState = 540)) or
								((vState = 572) and (hState = 560)) or
								((vState = 572) and (hState = 561)) or
								((vState = 572) and (hState = 565)) or
								((vState = 572) and (hState = 572)) or
								((vState = 572) and (hState = 579)) or
								((vState = 572) and (hState = 588)) or
								((vState = 572) and (hState = 589)) or
								((vState = 572) and (hState = 593)) or
								((vState = 573) and (hState = 524)) or
								((vState = 573) and (hState = 525)) or
								((vState = 573) and (hState = 526)) or
								((vState = 573) and (hState = 527)) or
								((vState = 573) and (hState = 562)) or
								((vState = 573) and (hState = 563)) or
								((vState = 573) and (hState = 564)) or
								((vState = 573) and (hState = 565)) or
								((vState = 573) and (hState = 573)) or
								((vState = 573) and (hState = 578)) or
								((vState = 573) and (hState = 587)) or
								((vState = 573) and (hState = 588)) or
								((vState = 573) and (hState = 589)) or
								((vState = 573) and (hState = 594)) or
								((vState = 574) and (hState = 523)) or
								((vState = 574) and (hState = 535)) or
								((vState = 574) and (hState = 562)) or
								((vState = 574) and (hState = 563)) or
								((vState = 574) and (hState = 564)) or
								((vState = 574) and (hState = 565)) or
								((vState = 574) and (hState = 566)) or
								((vState = 574) and (hState = 574)) or
								((vState = 574) and (hState = 577)) or
								((vState = 574) and (hState = 587)) or
								((vState = 574) and (hState = 588)) or
								((vState = 574) and (hState = 595)) or
								((vState = 575) and (hState = 511)) or
								((vState = 575) and (hState = 522)) or
								((vState = 575) and (hState = 535)) or
								((vState = 575) and (hState = 558)) or
								((vState = 575) and (hState = 562)) or
								((vState = 575) and (hState = 566)) or
								((vState = 575) and (hState = 567)) or
								((vState = 575) and (hState = 576)) or
								((vState = 575) and (hState = 577)) or
								((vState = 575) and (hState = 586)) or
								((vState = 575) and (hState = 587)) or
								((vState = 575) and (hState = 588)) or
								((vState = 576) and (hState = 510)) or
								((vState = 576) and (hState = 511)) or
								((vState = 576) and (hState = 512)) or
								((vState = 576) and (hState = 516)) or
								((vState = 576) and (hState = 517)) or
								((vState = 576) and (hState = 521)) or
								((vState = 576) and (hState = 522)) or
								((vState = 576) and (hState = 535)) or
								((vState = 576) and (hState = 558)) or
								((vState = 576) and (hState = 559)) or
								((vState = 576) and (hState = 567)) or
								((vState = 576) and (hState = 568)) or
								((vState = 576) and (hState = 576)) or
								((vState = 576) and (hState = 577)) or
								((vState = 576) and (hState = 585)) or
								((vState = 576) and (hState = 586)) or
								((vState = 576) and (hState = 587)) or
								((vState = 577) and (hState = 510)) or
								((vState = 577) and (hState = 511)) or
								((vState = 577) and (hState = 512)) or
								((vState = 577) and (hState = 513)) or
								((vState = 577) and (hState = 514)) or
								((vState = 577) and (hState = 515)) or
								((vState = 577) and (hState = 516)) or
								((vState = 577) and (hState = 517)) or
								((vState = 577) and (hState = 518)) or
								((vState = 577) and (hState = 519)) or
								((vState = 577) and (hState = 520)) or
								((vState = 577) and (hState = 521)) or
								((vState = 577) and (hState = 522)) or
								((vState = 577) and (hState = 531)) or
								((vState = 577) and (hState = 532)) or
								((vState = 577) and (hState = 533)) or
								((vState = 577) and (hState = 534)) or
								((vState = 577) and (hState = 535)) or
								((vState = 577) and (hState = 557)) or
								((vState = 577) and (hState = 558)) or
								((vState = 577) and (hState = 559)) or
								((vState = 577) and (hState = 567)) or
								((vState = 577) and (hState = 568)) or
								((vState = 577) and (hState = 576)) or
								((vState = 577) and (hState = 577)) or
								((vState = 577) and (hState = 584)) or
								((vState = 577) and (hState = 585)) or
								((vState = 577) and (hState = 586)) or
								((vState = 577) and (hState = 598)) or
								((vState = 578) and (hState = 515)) or
								((vState = 578) and (hState = 516)) or
								((vState = 578) and (hState = 517)) or
								((vState = 578) and (hState = 518)) or
								((vState = 578) and (hState = 519)) or
								((vState = 578) and (hState = 520)) or
								((vState = 578) and (hState = 521)) or
								((vState = 578) and (hState = 522)) or
								((vState = 578) and (hState = 531)) or
								((vState = 578) and (hState = 532)) or
								((vState = 578) and (hState = 533)) or
								((vState = 578) and (hState = 534)) or
								((vState = 578) and (hState = 535)) or
								((vState = 578) and (hState = 557)) or
								((vState = 578) and (hState = 558)) or
								((vState = 578) and (hState = 568)) or
								((vState = 578) and (hState = 569)) or
								((vState = 578) and (hState = 574)) or
								((vState = 578) and (hState = 578)) or
								((vState = 578) and (hState = 583)) or
								((vState = 578) and (hState = 584)) or
								((vState = 578) and (hState = 585)) or
								((vState = 578) and (hState = 586)) or
								((vState = 578) and (hState = 599)) or
								((vState = 579) and (hState = 516)) or
								((vState = 579) and (hState = 517)) or
								((vState = 579) and (hState = 525)) or
								((vState = 579) and (hState = 526)) or
								((vState = 579) and (hState = 527)) or
								((vState = 579) and (hState = 528)) or
								((vState = 579) and (hState = 529)) or
								((vState = 579) and (hState = 530)) or
								((vState = 579) and (hState = 531)) or
								((vState = 579) and (hState = 532)) or
								((vState = 579) and (hState = 533)) or
								((vState = 579) and (hState = 534)) or
								((vState = 579) and (hState = 535)) or
								((vState = 579) and (hState = 556)) or
								((vState = 579) and (hState = 557)) or
								((vState = 579) and (hState = 579)) or
								((vState = 579) and (hState = 583)) or
								((vState = 579) and (hState = 584)) or
								((vState = 579) and (hState = 585)) or
								((vState = 579) and (hState = 599)) or
								((vState = 580) and (hState = 517)) or
								((vState = 580) and (hState = 532)) or
								((vState = 580) and (hState = 533)) or
								((vState = 580) and (hState = 534)) or
								((vState = 580) and (hState = 535)) or
								((vState = 580) and (hState = 556)) or
								((vState = 580) and (hState = 583)) or
								((vState = 580) and (hState = 584)) or
								((vState = 580) and (hState = 585)) or
								((vState = 580) and (hState = 599)) or
								((vState = 581) and (hState = 517)) or
								((vState = 581) and (hState = 532)) or
								((vState = 581) and (hState = 533)) or
								((vState = 581) and (hState = 534)) or
								((vState = 581) and (hState = 535)) or
								((vState = 581) and (hState = 536)) or
								((vState = 581) and (hState = 537)) or
								((vState = 581) and (hState = 538)) or
								((vState = 581) and (hState = 572)) or
								((vState = 581) and (hState = 573)) or
								((vState = 581) and (hState = 581)) or
								((vState = 581) and (hState = 582)) or
								((vState = 581) and (hState = 583)) or
								((vState = 581) and (hState = 584)) or
								((vState = 581) and (hState = 599)) or
								((vState = 582) and (hState = 517)) or
								((vState = 582) and (hState = 532)) or
								((vState = 582) and (hState = 533)) or
								((vState = 582) and (hState = 534)) or
								((vState = 582) and (hState = 535)) or
								((vState = 582) and (hState = 536)) or
								((vState = 582) and (hState = 537)) or
								((vState = 582) and (hState = 538)) or
								((vState = 582) and (hState = 539)) or
								((vState = 582) and (hState = 540)) or
								((vState = 582) and (hState = 541)) or
								((vState = 582) and (hState = 542)) or
								((vState = 582) and (hState = 543)) or
								((vState = 582) and (hState = 544)) or
								((vState = 582) and (hState = 545)) or
								((vState = 582) and (hState = 572)) or
								((vState = 582) and (hState = 573)) or
								((vState = 582) and (hState = 581)) or
								((vState = 582) and (hState = 582)) or
								((vState = 582) and (hState = 583)) or
								((vState = 582) and (hState = 584)) or
								((vState = 582) and (hState = 599)) or
								((vState = 583) and (hState = 518)) or
								((vState = 583) and (hState = 534)) or
								((vState = 583) and (hState = 535)) or
								((vState = 583) and (hState = 536)) or
								((vState = 583) and (hState = 537)) or
								((vState = 583) and (hState = 538)) or
								((vState = 583) and (hState = 547)) or
								((vState = 583) and (hState = 548)) or
								((vState = 583) and (hState = 549)) or
								((vState = 583) and (hState = 550)) or
								((vState = 583) and (hState = 551)) or
								((vState = 583) and (hState = 552)) or
								((vState = 583) and (hState = 553)) or
								((vState = 583) and (hState = 554)) or
								((vState = 583) and (hState = 571)) or
								((vState = 583) and (hState = 572)) or
								((vState = 583) and (hState = 573)) or
								((vState = 583) and (hState = 574)) or
								((vState = 583) and (hState = 583)) or
								((vState = 583) and (hState = 584)) or
								((vState = 583) and (hState = 599)) or
								((vState = 584) and (hState = 519)) or
								((vState = 584) and (hState = 534)) or
								((vState = 584) and (hState = 535)) or
								((vState = 584) and (hState = 536)) or
								((vState = 584) and (hState = 537)) or
								((vState = 584) and (hState = 538)) or
								((vState = 584) and (hState = 550)) or
								((vState = 584) and (hState = 551)) or
								((vState = 584) and (hState = 574)) or
								((vState = 584) and (hState = 575)) or
								((vState = 584) and (hState = 579)) or
								((vState = 584) and (hState = 599)) or
								((vState = 585) and (hState = 535)) or
								((vState = 585) and (hState = 536)) or
								((vState = 585) and (hState = 574)) or
								((vState = 585) and (hState = 575)) or
								((vState = 585) and (hState = 576)) or
								((vState = 585) and (hState = 578)) or
								((vState = 585) and (hState = 579)) or
								((vState = 585) and (hState = 599)) or
								((vState = 586) and (hState = 536)) or
								((vState = 586) and (hState = 541)) or
								((vState = 586) and (hState = 576)) or
								((vState = 586) and (hState = 577)) or
								((vState = 586) and (hState = 578)) or
								((vState = 586) and (hState = 579)) or
								((vState = 587) and (hState = 536)) or
								((vState = 587) and (hState = 541)) or
								((vState = 587) and (hState = 548)) or
								((vState = 587) and (hState = 568)) or
								((vState = 587) and (hState = 576)) or
								((vState = 587) and (hState = 577)) or
								((vState = 587) and (hState = 578)) or
								((vState = 587) and (hState = 579)) or
								((vState = 588) and (hState = 536)) or
								((vState = 588) and (hState = 542)) or
								((vState = 588) and (hState = 547)) or
								((vState = 588) and (hState = 576)) or
								((vState = 588) and (hState = 577)) or
								((vState = 589) and (hState = 523)) or
								((vState = 589) and (hState = 537)) or
								((vState = 589) and (hState = 544)) or
								((vState = 589) and (hState = 545)) or
								((vState = 589) and (hState = 546)) or
								((vState = 589) and (hState = 567)) or
								((vState = 589) and (hState = 576)) or
								((vState = 589) and (hState = 577)) or
								((vState = 590) and (hState = 524)) or
								((vState = 590) and (hState = 537)) or
								((vState = 590) and (hState = 544)) or
								((vState = 590) and (hState = 545)) or
								((vState = 590) and (hState = 546)) or
								((vState = 590) and (hState = 578)) or
								((vState = 590) and (hState = 584)) or
								((vState = 591) and (hState = 525)) or
								((vState = 591) and (hState = 537)) or
								((vState = 591) and (hState = 538)) or
								((vState = 591) and (hState = 544)) or
								((vState = 591) and (hState = 545)) or
								((vState = 591) and (hState = 546)) or
								((vState = 591) and (hState = 574)) or
								((vState = 591) and (hState = 579)) or
								((vState = 591) and (hState = 585)) or
								((vState = 592) and (hState = 525)) or
								((vState = 592) and (hState = 526)) or
								((vState = 592) and (hState = 527)) or
								((vState = 592) and (hState = 537)) or
								((vState = 592) and (hState = 538)) or
								((vState = 592) and (hState = 539)) or
								((vState = 592) and (hState = 540)) or
								((vState = 592) and (hState = 541)) or
								((vState = 592) and (hState = 542)) or
								((vState = 592) and (hState = 543)) or
								((vState = 592) and (hState = 544)) or
								((vState = 592) and (hState = 545)) or
								((vState = 592) and (hState = 546)) or
								((vState = 592) and (hState = 547)) or
								((vState = 592) and (hState = 573)) or
								((vState = 592) and (hState = 574)) or
								((vState = 592) and (hState = 579)) or
								((vState = 592) and (hState = 585)) or
								((vState = 592) and (hState = 586)) or
								((vState = 593) and (hState = 527)) or
								((vState = 593) and (hState = 537)) or
								((vState = 593) and (hState = 538)) or
								((vState = 593) and (hState = 539)) or
								((vState = 593) and (hState = 540)) or
								((vState = 593) and (hState = 541)) or
								((vState = 593) and (hState = 547)) or
								((vState = 593) and (hState = 573)) or
								((vState = 594) and (hState = 537)) or
								((vState = 594) and (hState = 538)) or
								((vState = 594) and (hState = 539)) or
								((vState = 594) and (hState = 540)) or
								((vState = 594) and (hState = 541)) or
								((vState = 594) and (hState = 548)) or
								((vState = 594) and (hState = 563)) or
								((vState = 594) and (hState = 588)) or
								((vState = 595) and (hState = 537)) or
								((vState = 595) and (hState = 538)) or
								((vState = 595) and (hState = 539)) or
								((vState = 595) and (hState = 540)) or
								((vState = 595) and (hState = 541)) or
								((vState = 595) and (hState = 562)) or
								((vState = 595) and (hState = 572)) or
								((vState = 595) and (hState = 590)) or
								((vState = 596) and (hState = 529)) or
								((vState = 596) and (hState = 551)) or
								((vState = 596) and (hState = 583)) or
								((vState = 597) and (hState = 530)) or
								((vState = 597) and (hState = 542)) or
								((vState = 597) and (hState = 552)) or
								((vState = 597) and (hState = 583)) or
								((vState = 597) and (hState = 593)) or
								((vState = 598) and (hState = 530)) or
								((vState = 598) and (hState = 583)) or
								((vState = 598) and (hState = 593)) or
								((vState = 599) and (hState = 569)) or
								((vState = 599) and (hState = 583)) or
								((vState = 599) and (hState = 584)) or
								((vState = 600) and (hState = 532)) or
								((vState = 600) and (hState = 558)) or
								((vState = 600) and (hState = 569)) or
								((vState = 600) and (hState = 582)) or
								((vState = 600) and (hState = 583)) or
								((vState = 600) and (hState = 584)) or
								((vState = 600) and (hState = 585)) or
								((vState = 601) and (hState = 557)) or
								((vState = 601) and (hState = 558)) or
								((vState = 601) and (hState = 569)) or
								((vState = 601) and (hState = 582)) or
								((vState = 601) and (hState = 583)) or
								((vState = 602) and (hState = 546)) or
								((vState = 602) and (hState = 557)) or
								((vState = 602) and (hState = 558)) or
								((vState = 602) and (hState = 582)) or
								((vState = 602) and (hState = 583)) or
								((vState = 602) and (hState = 598)) or
								((vState = 603) and (hState = 546)) or
								((vState = 605) and (hState = 536)) or
								((vState = 605) and (hState = 547)) or
								((vState = 605) and (hState = 561)) or
								((vState = 605) and (hState = 572)) or
								((vState = 605) and (hState = 584)) or
								((vState = 606) and (hState = 537)) or
								((vState = 606) and (hState = 562)) or
								((vState = 606) and (hState = 584)) or
								((vState = 606) and (hState = 589)) or
								((vState = 607) and (hState = 553)) or
								((vState = 607) and (hState = 563)) or
								((vState = 607) and (hState = 573)) or
								((vState = 607) and (hState = 590)) or
								((vState = 608) and (hState = 553)) or
								((vState = 609) and (hState = 551)) or
								((vState = 609) and (hState = 585)) or
								((vState = 610) and (hState = 540)) or
								((vState = 610) and (hState = 551)) or
								((vState = 610) and (hState = 585)) or
								((vState = 610) and (hState = 595)) or
								((vState = 611) and (hState = 541)) or
								((vState = 611) and (hState = 551)) or
								((vState = 611) and (hState = 567)) or
								((vState = 611) and (hState = 579)) or
								((vState = 611) and (hState = 585)) or
								((vState = 611) and (hState = 593)) or
								((vState = 611) and (hState = 594)) or
								((vState = 611) and (hState = 595)) or
								((vState = 612) and (hState = 542)) or
								((vState = 612) and (hState = 550)) or
								((vState = 612) and (hState = 551)) or
								((vState = 612) and (hState = 552)) or
								((vState = 612) and (hState = 568)) or
								((vState = 612) and (hState = 579)) or
								((vState = 612) and (hState = 580)) or
								((vState = 612) and (hState = 594)) or
								((vState = 613) and (hState = 543)) or
								((vState = 613) and (hState = 549)) or
								((vState = 613) and (hState = 552)) or
								((vState = 613) and (hState = 568)) or
								((vState = 613) and (hState = 579)) or
								((vState = 613) and (hState = 580)) or
								((vState = 613) and (hState = 581)) or
								((vState = 613) and (hState = 594)) or
								((vState = 614) and (hState = 568)) or
								((vState = 614) and (hState = 579)) or
								((vState = 614) and (hState = 580)) or
								((vState = 614) and (hState = 581)) or
								((vState = 614) and (hState = 594)) or
								((vState = 615) and (hState = 568)) or
								((vState = 615) and (hState = 578)) or
								((vState = 615) and (hState = 579)) or
								((vState = 615) and (hState = 580)) or
								((vState = 615) and (hState = 581)) or
								((vState = 616) and (hState = 546)) or
								((vState = 616) and (hState = 547)) or
								((vState = 616) and (hState = 568)) or
								((vState = 616) and (hState = 578)) or
								((vState = 616) and (hState = 579)) or
								((vState = 616) and (hState = 580)) or
								((vState = 616) and (hState = 581)) or
								((vState = 616) and (hState = 593)) or
								((vState = 617) and (hState = 546)) or
								((vState = 617) and (hState = 547)) or
								((vState = 617) and (hState = 568)) or
								((vState = 617) and (hState = 578)) or
								((vState = 617) and (hState = 579)) or
								((vState = 617) and (hState = 580)) or
								((vState = 617) and (hState = 581)) or
								((vState = 617) and (hState = 588)) or
								((vState = 617) and (hState = 593)) or
								((vState = 617) and (hState = 597)) or
								((vState = 618) and (hState = 545)) or
								((vState = 618) and (hState = 546)) or
								((vState = 618) and (hState = 547)) or
								((vState = 618) and (hState = 556)) or
								((vState = 618) and (hState = 568)) or
								((vState = 618) and (hState = 578)) or
								((vState = 618) and (hState = 579)) or
								((vState = 618) and (hState = 580)) or
								((vState = 618) and (hState = 581)) or
								((vState = 618) and (hState = 588)) or
								((vState = 618) and (hState = 593)) or
								((vState = 618) and (hState = 594)) or
								((vState = 619) and (hState = 545)) or
								((vState = 619) and (hState = 546)) or
								((vState = 619) and (hState = 547)) or
								((vState = 619) and (hState = 578)) or
								((vState = 619) and (hState = 579)) or
								((vState = 619) and (hState = 580)) or
								((vState = 619) and (hState = 581)) or
								((vState = 619) and (hState = 588)) or
								((vState = 620) and (hState = 545)) or
								((vState = 620) and (hState = 546)) or
								((vState = 620) and (hState = 580)) or
								((vState = 620) and (hState = 581)) or
								((vState = 620) and (hState = 589)) or
								((vState = 620) and (hState = 590)) or
								((vState = 620) and (hState = 591)) or
								((vState = 621) and (hState = 544)) or
								((vState = 621) and (hState = 545)) or
								((vState = 621) and (hState = 546)) or
								((vState = 621) and (hState = 557)) or
								((vState = 621) and (hState = 567)) or
								((vState = 621) and (hState = 577)) or
								((vState = 621) and (hState = 581)) or
								((vState = 621) and (hState = 582)) or
								((vState = 621) and (hState = 583)) or
								((vState = 621) and (hState = 584)) or
								((vState = 621) and (hState = 585)) or
								((vState = 621) and (hState = 589)) or
								((vState = 621) and (hState = 590)) or
								((vState = 621) and (hState = 591)) or
								((vState = 622) and (hState = 542)) or
								((vState = 622) and (hState = 543)) or
								((vState = 622) and (hState = 544)) or
								((vState = 622) and (hState = 545)) or
								((vState = 622) and (hState = 546)) or
								((vState = 622) and (hState = 558)) or
								((vState = 622) and (hState = 567)) or
								((vState = 622) and (hState = 577)) or
								((vState = 622) and (hState = 581)) or
								((vState = 622) and (hState = 582)) or
								((vState = 622) and (hState = 583)) or
								((vState = 622) and (hState = 589)) or
								((vState = 622) and (hState = 590)) or
								((vState = 623) and (hState = 542)) or
								((vState = 623) and (hState = 543)) or
								((vState = 623) and (hState = 544)) or
								((vState = 623) and (hState = 545)) or
								((vState = 623) and (hState = 558)) or
								((vState = 623) and (hState = 567)) or
								((vState = 623) and (hState = 576)) or
								((vState = 623) and (hState = 577)) or
								((vState = 623) and (hState = 578)) or
								((vState = 623) and (hState = 582)) or
								((vState = 623) and (hState = 583)) or
								((vState = 623) and (hState = 589)) or
								((vState = 623) and (hState = 590)) or
								((vState = 624) and (hState = 542)) or
								((vState = 624) and (hState = 543)) or
								((vState = 624) and (hState = 544)) or
								((vState = 624) and (hState = 567)) or
								((vState = 624) and (hState = 576)) or
								((vState = 624) and (hState = 583)) or
								((vState = 624) and (hState = 589)) or
								((vState = 624) and (hState = 590)) or
								((vState = 625) and (hState = 541)) or
								((vState = 625) and (hState = 542)) or
								((vState = 625) and (hState = 543)) or
								((vState = 625) and (hState = 567)) or
								((vState = 625) and (hState = 573)) or
								((vState = 625) and (hState = 574)) or
								((vState = 625) and (hState = 575)) or
								((vState = 625) and (hState = 583)) or
								((vState = 625) and (hState = 589)) or
								((vState = 625) and (hState = 590)) or
								((vState = 626) and (hState = 540)) or
								((vState = 626) and (hState = 541)) or
								((vState = 626) and (hState = 542)) or
								((vState = 626) and (hState = 567)) or
								((vState = 626) and (hState = 573)) or
								((vState = 626) and (hState = 574)) or
								((vState = 626) and (hState = 575)) or
								((vState = 626) and (hState = 583)) or
								((vState = 626) and (hState = 589)) or
								((vState = 626) and (hState = 590)) or
								((vState = 627) and (hState = 539)) or
								((vState = 627) and (hState = 540)) or
								((vState = 627) and (hState = 541)) or
								((vState = 627) and (hState = 542)) or
								((vState = 627) and (hState = 561)) or
								((vState = 627) and (hState = 565)) or
								((vState = 627) and (hState = 573)) or
								((vState = 627) and (hState = 574)) or
								((vState = 627) and (hState = 575)) or
								((vState = 627) and (hState = 582)) or
								((vState = 627) and (hState = 583)) or
								((vState = 627) and (hState = 584)) or
								((vState = 627) and (hState = 590)) or
								((vState = 628) and (hState = 539)) or
								((vState = 628) and (hState = 540)) or
								((vState = 628) and (hState = 541)) or
								((vState = 628) and (hState = 560)) or
								((vState = 628) and (hState = 561)) or
								((vState = 628) and (hState = 562)) or
								((vState = 628) and (hState = 563)) or
								((vState = 628) and (hState = 564)) or
								((vState = 628) and (hState = 565)) or
								((vState = 628) and (hState = 573)) or
								((vState = 628) and (hState = 574)) or
								((vState = 628) and (hState = 575)) or
								((vState = 628) and (hState = 576)) or
								((vState = 628) and (hState = 577)) or
								((vState = 628) and (hState = 578)) or
								((vState = 628) and (hState = 583)) or
								((vState = 628) and (hState = 584)) or
								((vState = 628) and (hState = 590)) or
								((vState = 629) and (hState = 538)) or
								((vState = 629) and (hState = 539)) or
								((vState = 629) and (hState = 540)) or
								((vState = 629) and (hState = 566)) or
								((vState = 629) and (hState = 583)) or
								((vState = 629) and (hState = 584)) or
								((vState = 630) and (hState = 537)) or
								((vState = 630) and (hState = 538)) or
								((vState = 630) and (hState = 539)) or
								((vState = 630) and (hState = 566)) or
								((vState = 630) and (hState = 572)) or
								((vState = 630) and (hState = 584)) or
								((vState = 631) and (hState = 536)) or
								((vState = 631) and (hState = 537)) or
								((vState = 631) and (hState = 538)) or
								((vState = 631) and (hState = 570)) or
								((vState = 631) and (hState = 571)) or
								((vState = 631) and (hState = 572)) or
								((vState = 631) and (hState = 584)) or
								((vState = 631) and (hState = 585)) or
								((vState = 632) and (hState = 535)) or
								((vState = 632) and (hState = 536)) or
								((vState = 632) and (hState = 537)) or
								((vState = 632) and (hState = 538)) or
								((vState = 632) and (hState = 547)) or
								((vState = 632) and (hState = 548)) or
								((vState = 632) and (hState = 549)) or
								((vState = 632) and (hState = 571)) or
								((vState = 632) and (hState = 572)) or
								((vState = 632) and (hState = 573)) or
								((vState = 632) and (hState = 574)) or
								((vState = 632) and (hState = 575)) or
								((vState = 632) and (hState = 584)) or
								((vState = 632) and (hState = 585)) or
								((vState = 633) and (hState = 535)) or
								((vState = 633) and (hState = 536)) or
								((vState = 633) and (hState = 537)) or
								((vState = 633) and (hState = 547)) or
								((vState = 633) and (hState = 548)) or
								((vState = 633) and (hState = 577)) or
								((vState = 633) and (hState = 578)) or
								((vState = 633) and (hState = 579)) or
								((vState = 633) and (hState = 584)) or
								((vState = 633) and (hState = 585)) or
								((vState = 633) and (hState = 586)) or
								((vState = 634) and (hState = 534)) or
								((vState = 634) and (hState = 535)) or
								((vState = 634) and (hState = 536)) or
								((vState = 634) and (hState = 548)) or
								((vState = 634) and (hState = 569)) or
								((vState = 634) and (hState = 581)) or
								((vState = 634) and (hState = 582)) or
								((vState = 634) and (hState = 583)) or
								((vState = 634) and (hState = 584)) or
								((vState = 634) and (hState = 585)) or
								((vState = 634) and (hState = 586)) or
								((vState = 634) and (hState = 587)) or
								((vState = 634) and (hState = 588)) or
								((vState = 634) and (hState = 593)) or
								((vState = 635) and (hState = 534)) or
								((vState = 635) and (hState = 535)) or
								((vState = 635) and (hState = 536)) or
								((vState = 635) and (hState = 584)) or
								((vState = 635) and (hState = 585)) or
								((vState = 635) and (hState = 586)) or
								((vState = 635) and (hState = 587)) or
								((vState = 635) and (hState = 588)) or
								((vState = 635) and (hState = 593)) or
								((vState = 636) and (hState = 536)) or
								((vState = 636) and (hState = 584)) or
								((vState = 636) and (hState = 588)) or
								((vState = 636) and (hState = 593)) or
								((vState = 637) and (hState = 536)) or
								((vState = 637) and (hState = 552)) or
								((vState = 637) and (hState = 568)) or
								((vState = 637) and (hState = 584)) or
								((vState = 637) and (hState = 588)) or
								((vState = 637) and (hState = 589)) or
								((vState = 637) and (hState = 590)) or
								((vState = 637) and (hState = 591)) or
								((vState = 637) and (hState = 592)) or
								((vState = 637) and (hState = 593)) or
								((vState = 638) and (hState = 537)) or
								((vState = 638) and (hState = 553)) or
								((vState = 638) and (hState = 584)) or
								((vState = 638) and (hState = 589)) or
								((vState = 638) and (hState = 590)) or
								((vState = 638) and (hState = 591)) or
								((vState = 638) and (hState = 592)) or
								((vState = 638) and (hState = 593)) or
								((vState = 638) and (hState = 594)) or
								((vState = 639) and (hState = 540)) or
								((vState = 639) and (hState = 565)) or
								((vState = 639) and (hState = 566)) or
								((vState = 639) and (hState = 567)) or
								((vState = 639) and (hState = 584)) or
								((vState = 639) and (hState = 589)) or
								((vState = 639) and (hState = 590)) or
								((vState = 639) and (hState = 591)) or
								((vState = 639) and (hState = 592)) or
								((vState = 639) and (hState = 593)) or
								((vState = 639) and (hState = 594)) or
								((vState = 639) and (hState = 595)) or
								((vState = 639) and (hState = 596)) or
								((vState = 639) and (hState = 597)) or
								((vState = 640) and (hState = 565)) or
								((vState = 640) and (hState = 566)) or
								((vState = 640) and (hState = 589)) or
								((vState = 640) and (hState = 590)) or
								((vState = 640) and (hState = 591)) or
								((vState = 640) and (hState = 592)) or
								((vState = 640) and (hState = 593)) or
								((vState = 640) and (hState = 594)) or
								((vState = 640) and (hState = 595)) or
								((vState = 640) and (hState = 596)) or
								((vState = 640) and (hState = 597)) or
								((vState = 640) and (hState = 598)) or
								((vState = 641) and (hState = 565)) or
								((vState = 641) and (hState = 591)) or
								((vState = 641) and (hState = 592)) or
								((vState = 641) and (hState = 595)) or
								((vState = 642) and (hState = 557)) or
								((vState = 642) and (hState = 563)) or
								((vState = 642) and (hState = 564)) or
								((vState = 642) and (hState = 565)) or
								((vState = 642) and (hState = 585)) or
								((vState = 642) and (hState = 586)) or
								((vState = 642) and (hState = 595)) or
								((vState = 643) and (hState = 545)) or
								((vState = 643) and (hState = 563)) or
								((vState = 643) and (hState = 564)) or
								((vState = 643) and (hState = 585)) or
								((vState = 643) and (hState = 595)) or
								((vState = 644) and (hState = 547)) or
								((vState = 644) and (hState = 561)) or
								((vState = 644) and (hState = 562)) or
								((vState = 644) and (hState = 563)) or
								((vState = 644) and (hState = 564)) or
								((vState = 644) and (hState = 584)) or
								((vState = 644) and (hState = 585)) or
								((vState = 644) and (hState = 593)) or
								((vState = 644) and (hState = 594)) or
								((vState = 644) and (hState = 595)) or
								((vState = 645) and (hState = 562)) or
								((vState = 645) and (hState = 563)) or
								((vState = 645) and (hState = 585)) or
								((vState = 645) and (hState = 594)) or
								((vState = 645) and (hState = 595)) or
								((vState = 646) and (hState = 562)) or
								((vState = 646) and (hState = 563)) or
								((vState = 646) and (hState = 585)) or
								((vState = 646) and (hState = 594)) or
								((vState = 646) and (hState = 595)) or
								((vState = 647) and (hState = 563)) or
								((vState = 647) and (hState = 585)) or
								((vState = 647) and (hState = 595)) or
								((vState = 648) and (hState = 552)) or
								((vState = 648) and (hState = 563)) or
								((vState = 648) and (hState = 564)) or
								((vState = 648) and (hState = 579)) or
								((vState = 648) and (hState = 585)) or
								((vState = 648) and (hState = 595)) or
								((vState = 648) and (hState = 596)) or
								((vState = 649) and (hState = 553)) or
								((vState = 649) and (hState = 554)) or
								((vState = 649) and (hState = 577)) or
								((vState = 649) and (hState = 595)) or
								((vState = 649) and (hState = 596)) or
								((vState = 650) and (hState = 577)) or
								((vState = 654) and (hState = 572)) or
								((vState = 655) and (hState = 563)) or
								((vState = 655) and (hState = 573)) or
								((vState = 655) and (hState = 584)) or
								((vState = 655) and (hState = 585)) or
								((vState = 655) and (hState = 586)) or
								((vState = 656) and (hState = 585)) or
								((vState = 656) and (hState = 586)) or
								((vState = 658) and (hState = 567)) or
								((vState = 659) and (hState = 568)) or
								((vState = 659) and (hState = 578)) or
								((vState = 659) and (hState = 588)) or
								((vState = 659) and (hState = 589)) or
								((vState = 660) and (hState = 579)) or
								((vState = 660) and (hState = 588)) or
								((vState = 660) and (hState = 589)) or
								((vState = 660) and (hState = 590)) or
								((vState = 661) and (hState = 588)) or
								((vState = 662) and (hState = 588)) or
								((vState = 663) and (hState = 588)) or
								((vState = 663) and (hState = 594)) or
								((vState = 664) and (hState = 583)) or
								((vState = 664) and (hState = 588)) or
								((vState = 664) and (hState = 595)) or
								((vState = 665) and (hState = 585)) or
								((vState = 665) and (hState = 586)) or
								((vState = 665) and (hState = 587)) or
								((vState = 665) and (hState = 588)) or
								((vState = 666) and (hState = 587)) or
								((vState = 666) and (hState = 588)) or
								((vState = 667) and (hState = 588)) else (others => '0');
end architecture me;
